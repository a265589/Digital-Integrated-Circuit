.SUBCKT Accumulator VSS VDD  clk rst_n in_valid partial_sum[12] partial_sum[11] partial_sum[10] partial_sum[9] partial_sum[8] partial_sum[7] partial_sum[6] partial_sum[5] partial_sum[4] partial_sum[3] partial_sum[2] partial_sum[1] partial_sum[0] result[12] result[11] result[10] result[9] result[8] result[7] result[6] result[5] result[4] result[3] result[2] result[1] result[0]
Xresult_reg_12_ VSS VDD  clk N_30  n2 n30 n14 ASYNC_DFFHx1_ASAP7_75t_R
Xresult_reg_11_ VSS VDD  clk N_29  n2 n56 n13 ASYNC_DFFHx1_ASAP7_75t_R
Xresult_reg_10_ VSS VDD  clk N_28  n2 n28 n12 ASYNC_DFFHx1_ASAP7_75t_R
Xresult_reg_9_ VSS VDD   clk N_27  n2 n57 n11 ASYNC_DFFHx1_ASAP7_75t_R
Xresult_reg_8_ VSS VDD   clk N_26  n2 n29 n10 ASYNC_DFFHx1_ASAP7_75t_R
Xresult_reg_7_ VSS VDD   clk N_25  n2 n25 n9 ASYNC_DFFHx1_ASAP7_75t_R
Xresult_reg_6_ VSS VDD   clk N_24  n2 n55 n8 ASYNC_DFFHx1_ASAP7_75t_R
Xresult_reg_5_ VSS VDD   clk N_23  n2 n27 n7 ASYNC_DFFHx1_ASAP7_75t_R
Xresult_reg_4_ VSS VDD   clk N_22  n2 n32 n6 ASYNC_DFFHx1_ASAP7_75t_R
Xresult_reg_3_ VSS VDD   clk N_21  n2 n54 n5 ASYNC_DFFHx1_ASAP7_75t_R
Xresult_reg_2_ VSS VDD   clk N_20  n2 n15 n4 ASYNC_DFFHx1_ASAP7_75t_R
Xresult_reg_1_ VSS VDD   clk N_19  n2 n31 n3 ASYNC_DFFHx1_ASAP7_75t_R
Xresult_reg_0_ VSS VDD   clk N_18  n2 n26 n1 ASYNC_DFFHx1_ASAP7_75t_R
XU31 VSS VDD  n37 result[7] INVx1_ASAP7_75t_R
XU32 VSS VDD  n36 result[5] INVx1_ASAP7_75t_R
XU33 VSS VDD  n35 result[3] INVx1_ASAP7_75t_R
XU34 VSS VDD  n38 result[9] INVx1_ASAP7_75t_R
XU35 VSS VDD  n116 result[10] INVx3_ASAP7_75t_R
XU36 VSS VDD  n40 result[1] INVx1_ASAP7_75t_R
XU37 VSS VDD  n117 result[8] INVx3_ASAP7_75t_R
XU38 VSS VDD  n118 result[6] INVx3_ASAP7_75t_R
XU39 VSS VDD  n119 result[4] INVx3_ASAP7_75t_R
XU40 VSS VDD  n120 result[2] INVx3_ASAP7_75t_R
XU41 VSS VDD  n121 result[0] INVx2_ASAP7_75t_R
XU42 VSS VDD  n1 n121 BUFx3_ASAP7_75t_R
XU43 VSS VDD  n11 n38 BUFx5_ASAP7_75t_R
XU44 VSS VDD  n3 n40 BUFx5_ASAP7_75t_R
XU45 VSS VDD  n5 n35 BUFx5_ASAP7_75t_R
XU46 VSS VDD  n7 n36 BUFx5_ASAP7_75t_R
XU47 VSS VDD  n9 n37 BUFx5_ASAP7_75t_R
XU48 VSS VDD  in_valid n16 INVx8_ASAP7_75t_R
XU49 VSS VDD  in_valid n17 INVx8_ASAP7_75t_R
XU50 VSS VDD  in_valid n18 INVx8_ASAP7_75t_R
XU51 VSS VDD  in_valid n19 INVx8_ASAP7_75t_R
XU52 VSS VDD  in_valid n20 INVx8_ASAP7_75t_R
XU53 VSS VDD  result[0] partial_sum[1] n21 NAND2xp33_ASAP7_75t_R
XU54 VSS VDD  in_valid n22 INVx8_ASAP7_75t_R
XU55 VSS VDD  in_valid n23 INVx8_ASAP7_75t_R
XU56 VSS VDD  result[0] partial_sum[1] n24 AND2x2_ASAP7_75t_R
XU57 VSS VDD  rst_n n25 INVx8_ASAP7_75t_R
XU58 VSS VDD  rst_n n26 INVx8_ASAP7_75t_R
XU59 VSS VDD  rst_n n27 INVx8_ASAP7_75t_R
XU60 VSS VDD  rst_n n28 INVx8_ASAP7_75t_R
XU61 VSS VDD  rst_n n29 INVx8_ASAP7_75t_R
XU62 VSS VDD  rst_n n30 INVx8_ASAP7_75t_R
XU63 VSS VDD  rst_n n31 INVx8_ASAP7_75t_R
XU64 VSS VDD  rst_n n32 INVx8_ASAP7_75t_R
XU65 VSS VDD  n6 n119 BUFx5_ASAP7_75t_R
XU66 VSS VDD  n10 n117 BUFx5_ASAP7_75t_R
XU67 VSS VDD  n12 n116 BUFx5_ASAP7_75t_R
XU68 VSS VDD  n13 n33 BUFx3_ASAP7_75t_R
XU69 VSS VDD  n8 n118 BUFx5_ASAP7_75t_R
XU70 VSS VDD  n4 n120 BUFx5_ASAP7_75t_R
XU71 VSS VDD  partial_sum[10] n45 INVx8_ASAP7_75t_R
XU72 VSS VDD  partial_sum[10] n106 INVx8_ASAP7_75t_R
XU73 VSS VDD  partial_sum[8] n46 INVx8_ASAP7_75t_R
XU74 VSS VDD  partial_sum[8] n95 INVx8_ASAP7_75t_R
XU75 VSS VDD  partial_sum[6] n47 INVx8_ASAP7_75t_R
XU76 VSS VDD  partial_sum[6] n84 INVx8_ASAP7_75t_R
XU77 VSS VDD  partial_sum[4] n48 INVx8_ASAP7_75t_R
XU78 VSS VDD  partial_sum[4] n73 INVx8_ASAP7_75t_R
XU79 VSS VDD  partial_sum[2] n49 INVx8_ASAP7_75t_R
XU80 VSS VDD  partial_sum[2] n63 INVx8_ASAP7_75t_R
XU81 VSS VDD  in_valid n50 INVx8_ASAP7_75t_R
XU82 VSS VDD  in_valid n51 INVx8_ASAP7_75t_R
XU83 VSS VDD  in_valid n52 INVx8_ASAP7_75t_R
XU84 VSS VDD  in_valid n53 INVx8_ASAP7_75t_R
XU85 VSS VDD  in_valid n115 INVx8_ASAP7_75t_R
XU86 VSS VDD  rst_n n54 INVx8_ASAP7_75t_R
XU87 VSS VDD  rst_n n55 INVx8_ASAP7_75t_R
XU88 VSS VDD  rst_n n56 INVx8_ASAP7_75t_R
XU89 VSS VDD  rst_n n57 INVx8_ASAP7_75t_R
XU90 VSS VDD  rst_n n15 INVx8_ASAP7_75t_R
XU91 VSS VDD  n2 TIELOx1_ASAP7_75t_R
XU92 VSS VDD  n14 result[12] INVxp33_ASAP7_75t_R
XU93 VSS VDD  n33 result[11] INVxp33_ASAP7_75t_R
XU94 VSS VDD  in_valid partial_sum[0] N_18 AND2x2_ASAP7_75t_R
XU95 VSS VDD  result[0] partial_sum[1] n58 NOR2xp33_ASAP7_75t_R
XU96 VSS VDD  n58 n22 n24 N_19 NOR3xp33_ASAP7_75t_R
XU97 VSS VDD  result[1] partial_sum[2] n60 NOR2xp33_ASAP7_75t_R
XU98 VSS VDD  n40 n63 n59 NOR2xp33_ASAP7_75t_R
XU99 VSS VDD  n60 n59 n61 NOR2xp33_ASAP7_75t_R
XU100 VSS VDD  n61 n24 A0  n62 HAxp5_ASAP7_75t_R
XU101 VSS VDD  n16 n62 N_20 NOR2xp33_ASAP7_75t_R
XU102 VSS VDD  n40 n21 n49 n68 MAJIxp5_ASAP7_75t_R
XU103 VSS VDD  result[2] partial_sum[3] n65 AND2x2_ASAP7_75t_R
XU104 VSS VDD  result[2] partial_sum[3] n64 NOR2xp33_ASAP7_75t_R
XU105 VSS VDD  n65 n64 n66 NOR2xp33_ASAP7_75t_R
XU106 VSS VDD  n68 n66 A1  n67 HAxp5_ASAP7_75t_R
XU107 VSS VDD  n50 n67 N_21 NOR2xp33_ASAP7_75t_R
XU108 VSS VDD  result[2] partial_sum[3] n68 n74 MAJIxp5_ASAP7_75t_R
XU109 VSS VDD  n35 n73 n70 NOR2xp33_ASAP7_75t_R
XU110 VSS VDD  result[3] partial_sum[4] n69 NOR2xp33_ASAP7_75t_R
XU111 VSS VDD  n70 n69 n71 NOR2xp33_ASAP7_75t_R
XU112 VSS VDD  n74 n71 n72 XOR2xp5_ASAP7_75t_R
XU113 VSS VDD  n115 n72 N_22 NOR2xp33_ASAP7_75t_R
XU114 VSS VDD  n35 n74 n48 n79 MAJIxp5_ASAP7_75t_R
XU115 VSS VDD  result[4] partial_sum[5] n76 AND2x2_ASAP7_75t_R
XU116 VSS VDD  result[4] partial_sum[5] n75 NOR2xp33_ASAP7_75t_R
XU117 VSS VDD  n76 n75 n77 NOR2xp33_ASAP7_75t_R
XU118 VSS VDD  n79 n77 A2  n78 HAxp5_ASAP7_75t_R
XU119 VSS VDD  n23 n78 N_23 NOR2xp33_ASAP7_75t_R
XU120 VSS VDD  result[4] partial_sum[5] n79 n85 MAJIxp5_ASAP7_75t_R
XU121 VSS VDD  n36 n84 n81 NOR2xp33_ASAP7_75t_R
XU122 VSS VDD  result[5] partial_sum[6] n80 NOR2xp33_ASAP7_75t_R
XU123 VSS VDD  n81 n80 n82 NOR2xp33_ASAP7_75t_R
XU124 VSS VDD  n85 n82 n83 XOR2xp5_ASAP7_75t_R
XU125 VSS VDD  n51 n83 N_24 NOR2xp33_ASAP7_75t_R
XU126 VSS VDD  n36 n85 n47 n90 MAJIxp5_ASAP7_75t_R
XU127 VSS VDD  result[6] partial_sum[7] n87 AND2x2_ASAP7_75t_R
XU128 VSS VDD  result[6] partial_sum[7] n86 NOR2xp33_ASAP7_75t_R
XU129 VSS VDD  n87 n86 n88 NOR2xp33_ASAP7_75t_R
XU130 VSS VDD  n90 n88 A3  n89 HAxp5_ASAP7_75t_R
XU131 VSS VDD  n17 n89 N_25 NOR2xp33_ASAP7_75t_R
XU132 VSS VDD  result[6] partial_sum[7] n90 n96 MAJIxp5_ASAP7_75t_R
XU133 VSS VDD  n37 n95 n92 NOR2xp33_ASAP7_75t_R
XU134 VSS VDD  result[7] partial_sum[8] n91 NOR2xp33_ASAP7_75t_R
XU135 VSS VDD  n92 n91 n93 NOR2xp33_ASAP7_75t_R
XU136 VSS VDD  n96 n93 n94 XOR2xp5_ASAP7_75t_R
XU137 VSS VDD  n20 n94 N_26 NOR2xp33_ASAP7_75t_R
XU138 VSS VDD  n37 n96 n46 n101 MAJIxp5_ASAP7_75t_R
XU139 VSS VDD  result[8] partial_sum[9] n98 AND2x2_ASAP7_75t_R
XU140 VSS VDD  result[8] partial_sum[9] n97 NOR2xp33_ASAP7_75t_R
XU141 VSS VDD  n98 n97 n99 NOR2xp33_ASAP7_75t_R
XU142 VSS VDD  n101 n99 A4  n100 HAxp5_ASAP7_75t_R
XU143 VSS VDD  n18 n100 N_27 NOR2xp33_ASAP7_75t_R
XU144 VSS VDD  result[8] partial_sum[9] n101 n107 MAJIxp5_ASAP7_75t_R
XU145 VSS VDD  n38 n106 n103 NOR2xp33_ASAP7_75t_R
XU146 VSS VDD  result[9] partial_sum[10] n102 NOR2xp33_ASAP7_75t_R
XU147 VSS VDD  n103 n102 n104 NOR2xp33_ASAP7_75t_R
XU148 VSS VDD  n107 n104 n105 XOR2xp5_ASAP7_75t_R
XU149 VSS VDD  n53 n105 N_28 NOR2xp33_ASAP7_75t_R
XU150 VSS VDD  n38 n107 n45 n112 MAJIxp5_ASAP7_75t_R
XU151 VSS VDD  result[10] partial_sum[11] n109 NOR2xp33_ASAP7_75t_R
XU152 VSS VDD  result[10] partial_sum[11] n108 AND2x2_ASAP7_75t_R
XU153 VSS VDD  n109 n108 n110 NOR2xp33_ASAP7_75t_R
XU154 VSS VDD  n112 n110 A5  n111 HAxp5_ASAP7_75t_R
XU155 VSS VDD  n19 n111 N_29 NOR2xp33_ASAP7_75t_R
XU156 VSS VDD  result[10] partial_sum[11] n112 n113 MAJIxp5_ASAP7_75t_R
XU157 VSS VDD  partial_sum[12] n113 n33 A6  n114 FAx1_ASAP7_75t_R
XU158 VSS VDD  n52 n114 N_30 NOR2xp33_ASAP7_75t_R
.ENDS


