.SUBCKT Adder_tree VSS VDD  in[127] in[126] in[125] in[124] in[123] in[122] in[121] in[120] in[119] in[118] in[117] in[116] in[115] in[114] in[113] in[112] in[111] in[110] in[109] in[108] in[107] in[106] in[105] in[104] in[103] in[102] in[101] in[100] in[99] in[98] in[97] in[96] in[95] in[94] in[93] in[92] in[91] in[90] in[89] in[88] in[87] in[86] in[85] in[84] in[83] in[82] in[81] in[80] in[79] in[78] in[77] in[76] in[75] in[74] in[73] in[72] in[71] in[70] in[69] in[68] in[67] in[66] in[65] in[64] in[63] in[62] in[61] in[60] in[59] in[58] in[57] in[56] in[55] in[54] in[53] in[52] in[51] in[50] in[49] in[48] in[47] in[46] in[45] in[44] in[43] in[42] in[41] in[40] in[39] in[38] in[37] in[36] in[35] in[34] in[33] in[32] in[31] in[30] in[29] in[28] in[27] in[26] in[25] in[24] in[23] in[22] in[21] in[20] in[19] in[18] in[17] in[16] in[15] in[14] in[13] in[12] in[11] in[10] in[9] in[8] in[7] in[6] in[5] in[4] in[3] in[2] in[1] in[0] out[12] out[11] out[10] out[9] out[8] out[7] out[6] out[5] out[4] out[3] out[2] out[1] out[0]
XDP_OP_94J1_122_9915_U198 VSS VDD  in[4] in[28] in[36] DP_OP_94J1_122_9915_n299 DP_OP_94J1_122_9915_n300 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U197 VSS VDD  in[44] in[52] in[60] DP_OP_94J1_122_9915_n297 DP_OP_94J1_122_9915_n298 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U196 VSS VDD  in[68] in[76] in[84] DP_OP_94J1_122_9915_n295 DP_OP_94J1_122_9915_n296 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U195 VSS VDD  in[92] in[100] in[108] DP_OP_94J1_122_9915_n293 DP_OP_94J1_122_9915_n294 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U194 VSS VDD  in[116] in[124] in[120] DP_OP_94J1_122_9915_n291 DP_OP_94J1_122_9915_n292 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U193 VSS VDD  in[112] in[104] in[96] DP_OP_94J1_122_9915_n289 DP_OP_94J1_122_9915_n290 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U192 VSS VDD  in[88] in[80] in[72] DP_OP_94J1_122_9915_n287 DP_OP_94J1_122_9915_n288 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U191 VSS VDD  in[64] in[56] in[48] DP_OP_94J1_122_9915_n285 DP_OP_94J1_122_9915_n286 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U190 VSS VDD  in[40] in[0] in[32] DP_OP_94J1_122_9915_n283 DP_OP_94J1_122_9915_n284 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U189 VSS VDD  in[24] in[8] in[16] DP_OP_94J1_122_9915_n281 DP_OP_94J1_122_9915_n282 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U187 VSS VDD  DP_OP_94J1_122_9915_n284 DP_OP_94J1_122_9915_n278 DP_OP_94J1_122_9915_n286 DP_OP_94J1_122_9915_n279 DP_OP_94J1_122_9915_n280 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U186 VSS VDD  DP_OP_94J1_122_9915_n282 DP_OP_94J1_122_9915_n288 DP_OP_94J1_122_9915_n290 DP_OP_94J1_122_9915_n276 DP_OP_94J1_122_9915_n277 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U185 VSS VDD  DP_OP_94J1_122_9915_n292 DP_OP_94J1_122_9915_n294 DP_OP_94J1_122_9915_n296 DP_OP_94J1_122_9915_n274 DP_OP_94J1_122_9915_n275 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U183 VSS VDD  DP_OP_94J1_122_9915_n298 DP_OP_94J1_122_9915_n300 DP_OP_94J1_122_9915_n271 DP_OP_94J1_122_9915_n272 DP_OP_94J1_122_9915_n273 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U180 VSS VDD  in[21] in[29] in[37] DP_OP_94J1_122_9915_n267 DP_OP_94J1_122_9915_n268 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U179 VSS VDD  in[45] in[53] in[61] DP_OP_94J1_122_9915_n265 DP_OP_94J1_122_9915_n266 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U178 VSS VDD  in[69] in[77] in[85] DP_OP_94J1_122_9915_n263 DP_OP_94J1_122_9915_n264 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U177 VSS VDD  in[93] in[101] in[109] DP_OP_94J1_122_9915_n261 DP_OP_94J1_122_9915_n262 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U176 VSS VDD  in[117] in[81] in[1] DP_OP_94J1_122_9915_n259 DP_OP_94J1_122_9915_n260 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U175 VSS VDD  in[125] in[89] in[121] DP_OP_94J1_122_9915_n257 DP_OP_94J1_122_9915_n258 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U174 VSS VDD  in[9] in[65] in[17] DP_OP_94J1_122_9915_n255 DP_OP_94J1_122_9915_n256 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U173 VSS VDD  in[113] in[97] in[25] DP_OP_94J1_122_9915_n253 DP_OP_94J1_122_9915_n254 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U172 VSS VDD  in[105] in[33] in[73] DP_OP_94J1_122_9915_n251 DP_OP_94J1_122_9915_n252 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U171 VSS VDD  in[57] in[41] in[49] DP_OP_94J1_122_9915_n249 DP_OP_94J1_122_9915_n250 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U169 VSS VDD  DP_OP_94J1_122_9915_n299 DP_OP_94J1_122_9915_n246 DP_OP_94J1_122_9915_n297 DP_OP_94J1_122_9915_n247 DP_OP_94J1_122_9915_n248 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U167 VSS VDD  DP_OP_94J1_122_9915_n295 DP_OP_94J1_122_9915_n283 DP_OP_94J1_122_9915_n243 DP_OP_94J1_122_9915_n244 DP_OP_94J1_122_9915_n245 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U166 VSS VDD  DP_OP_94J1_122_9915_n285 DP_OP_94J1_122_9915_n281 DP_OP_94J1_122_9915_n287 DP_OP_94J1_122_9915_n241 DP_OP_94J1_122_9915_n242 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U165 VSS VDD  DP_OP_94J1_122_9915_n289 DP_OP_94J1_122_9915_n291 DP_OP_94J1_122_9915_n293 DP_OP_94J1_122_9915_n239 DP_OP_94J1_122_9915_n240 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U164 VSS VDD  DP_OP_94J1_122_9915_n260 DP_OP_94J1_122_9915_n250 DP_OP_94J1_122_9915_n262 DP_OP_94J1_122_9915_n237 DP_OP_94J1_122_9915_n238 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U163 VSS VDD  DP_OP_94J1_122_9915_n258 DP_OP_94J1_122_9915_n252 DP_OP_94J1_122_9915_n256 DP_OP_94J1_122_9915_n235 DP_OP_94J1_122_9915_n236 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U162 VSS VDD  DP_OP_94J1_122_9915_n266 DP_OP_94J1_122_9915_n254 DP_OP_94J1_122_9915_n264 DP_OP_94J1_122_9915_n233 DP_OP_94J1_122_9915_n234 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U160 VSS VDD  DP_OP_94J1_122_9915_n279 DP_OP_94J1_122_9915_n248 DP_OP_94J1_122_9915_n230 DP_OP_94J1_122_9915_n231 DP_OP_94J1_122_9915_n232 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U159 VSS VDD  DP_OP_94J1_122_9915_n240 DP_OP_94J1_122_9915_n242 DP_OP_94J1_122_9915_n245 DP_OP_94J1_122_9915_n228 DP_OP_94J1_122_9915_n229 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U158 VSS VDD  DP_OP_94J1_122_9915_n274 DP_OP_94J1_122_9915_n276 DP_OP_94J1_122_9915_n238 DP_OP_94J1_122_9915_n226 DP_OP_94J1_122_9915_n227 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U156 VSS VDD  DP_OP_94J1_122_9915_n234 DP_OP_94J1_122_9915_n236 DP_OP_94J1_122_9915_n223 DP_OP_94J1_122_9915_n224 DP_OP_94J1_122_9915_n225 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U154 VSS VDD  DP_OP_94J1_122_9915_n227 DP_OP_94J1_122_9915_n229 DP_OP_94J1_122_9915_n220 DP_OP_94J1_122_9915_n221 DP_OP_94J1_122_9915_n222 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U150 VSS VDD  in[22] in[30] in[38] DP_OP_94J1_122_9915_n215 DP_OP_94J1_122_9915_n216 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U149 VSS VDD  in[46] in[54] in[62] DP_OP_94J1_122_9915_n213 DP_OP_94J1_122_9915_n214 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U148 VSS VDD  in[2] in[106] in[10] DP_OP_94J1_122_9915_n211 DP_OP_94J1_122_9915_n212 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U147 VSS VDD  in[70] in[18] in[78] DP_OP_94J1_122_9915_n209 DP_OP_94J1_122_9915_n210 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U146 VSS VDD  in[86] in[26] in[34] DP_OP_94J1_122_9915_n207 DP_OP_94J1_122_9915_n208 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U145 VSS VDD  in[94] in[122] in[102] DP_OP_94J1_122_9915_n205 DP_OP_94J1_122_9915_n206 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U144 VSS VDD  in[110] in[42] in[118] DP_OP_94J1_122_9915_n203 DP_OP_94J1_122_9915_n204 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U143 VSS VDD  in[126] in[50] in[114] DP_OP_94J1_122_9915_n201 DP_OP_94J1_122_9915_n202 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U142 VSS VDD  in[58] in[90] in[66] DP_OP_94J1_122_9915_n199 DP_OP_94J1_122_9915_n200 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U141 VSS VDD  in[98] in[74] in[82] DP_OP_94J1_122_9915_n197 DP_OP_94J1_122_9915_n198 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U139 VSS VDD  DP_OP_94J1_122_9915_n267 DP_OP_94J1_122_9915_n194 DP_OP_94J1_122_9915_n265 DP_OP_94J1_122_9915_n195 DP_OP_94J1_122_9915_n196 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U137 VSS VDD  DP_OP_94J1_122_9915_n263 DP_OP_94J1_122_9915_n249 DP_OP_94J1_122_9915_n191 DP_OP_94J1_122_9915_n192 DP_OP_94J1_122_9915_n193 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U136 VSS VDD  DP_OP_94J1_122_9915_n261 DP_OP_94J1_122_9915_n257 DP_OP_94J1_122_9915_n251 DP_OP_94J1_122_9915_n189 DP_OP_94J1_122_9915_n190 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U135 VSS VDD  DP_OP_94J1_122_9915_n259 DP_OP_94J1_122_9915_n253 DP_OP_94J1_122_9915_n255 DP_OP_94J1_122_9915_n187 DP_OP_94J1_122_9915_n188 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U133 VSS VDD  DP_OP_94J1_122_9915_n241 DP_OP_94J1_122_9915_n247 DP_OP_94J1_122_9915_n184 DP_OP_94J1_122_9915_n185 DP_OP_94J1_122_9915_n186 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U131 VSS VDD  DP_OP_94J1_122_9915_n210 DP_OP_94J1_122_9915_n202 DP_OP_94J1_122_9915_n181 DP_OP_94J1_122_9915_n182 DP_OP_94J1_122_9915_n183 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U130 VSS VDD  DP_OP_94J1_122_9915_n214 DP_OP_94J1_122_9915_n204 DP_OP_94J1_122_9915_n216 DP_OP_94J1_122_9915_n179 DP_OP_94J1_122_9915_n180 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U129 VSS VDD  DP_OP_94J1_122_9915_n212 DP_OP_94J1_122_9915_n200 DP_OP_94J1_122_9915_n206 DP_OP_94J1_122_9915_n177 DP_OP_94J1_122_9915_n178 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U127 VSS VDD  DP_OP_94J1_122_9915_n244 DP_OP_94J1_122_9915_n196 DP_OP_94J1_122_9915_n174 DP_OP_94J1_122_9915_n175 DP_OP_94J1_122_9915_n176 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U126 VSS VDD  DP_OP_94J1_122_9915_n190 DP_OP_94J1_122_9915_n188 DP_OP_94J1_122_9915_n193 DP_OP_94J1_122_9915_n172 DP_OP_94J1_122_9915_n173 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U125 VSS VDD  DP_OP_94J1_122_9915_n233 DP_OP_94J1_122_9915_n237 DP_OP_94J1_122_9915_n235 DP_OP_94J1_122_9915_n170 DP_OP_94J1_122_9915_n171 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U123 VSS VDD  DP_OP_94J1_122_9915_n228 DP_OP_94J1_122_9915_n231 DP_OP_94J1_122_9915_n167 DP_OP_94J1_122_9915_n168 DP_OP_94J1_122_9915_n169 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U121 VSS VDD  DP_OP_94J1_122_9915_n180 DP_OP_94J1_122_9915_n178 DP_OP_94J1_122_9915_n164 DP_OP_94J1_122_9915_n165 DP_OP_94J1_122_9915_n166 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U120 VSS VDD  DP_OP_94J1_122_9915_n226 DP_OP_94J1_122_9915_n176 DP_OP_94J1_122_9915_n171 DP_OP_94J1_122_9915_n162 DP_OP_94J1_122_9915_n163 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U119 VSS VDD  DP_OP_94J1_122_9915_n224 DP_OP_94J1_122_9915_n173 DP_OP_94J1_122_9915_n166 DP_OP_94J1_122_9915_n160 DP_OP_94J1_122_9915_n161 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U118 VSS VDD  DP_OP_94J1_122_9915_n221 DP_OP_94J1_122_9915_n169 DP_OP_94J1_122_9915_n163 DP_OP_94J1_122_9915_n158 DP_OP_94J1_122_9915_n159 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U114 VSS VDD  in[23] in[31] in[39] DP_OP_94J1_122_9915_n153 DP_OP_94J1_122_9915_n154 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U113 VSS VDD  in[47] in[115] in[55] DP_OP_94J1_122_9915_n151 DP_OP_94J1_122_9915_n152 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U112 VSS VDD  in[63] in[3] in[71] DP_OP_94J1_122_9915_n149 DP_OP_94J1_122_9915_n150 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U111 VSS VDD  in[79] in[99] in[11] DP_OP_94J1_122_9915_n147 DP_OP_94J1_122_9915_n148 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U110 VSS VDD  in[19] in[107] in[87] DP_OP_94J1_122_9915_n145 DP_OP_94J1_122_9915_n146 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U109 VSS VDD  in[95] in[27] in[103] DP_OP_94J1_122_9915_n143 DP_OP_94J1_122_9915_n144 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U108 VSS VDD  in[111] in[35] in[119] DP_OP_94J1_122_9915_n141 DP_OP_94J1_122_9915_n142 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U107 VSS VDD  in[127] in[43] in[123] DP_OP_94J1_122_9915_n139 DP_OP_94J1_122_9915_n140 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U106 VSS VDD  in[91] in[51] in[83] DP_OP_94J1_122_9915_n137 DP_OP_94J1_122_9915_n138 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U105 VSS VDD  in[75] in[59] in[67] DP_OP_94J1_122_9915_n135 DP_OP_94J1_122_9915_n136 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U103 VSS VDD  DP_OP_94J1_122_9915_n215 DP_OP_94J1_122_9915_n132 DP_OP_94J1_122_9915_n213 DP_OP_94J1_122_9915_n133 DP_OP_94J1_122_9915_n134 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U101 VSS VDD  DP_OP_94J1_122_9915_n211 DP_OP_94J1_122_9915_n197 DP_OP_94J1_122_9915_n129 DP_OP_94J1_122_9915_n130 DP_OP_94J1_122_9915_n131 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U100 VSS VDD  DP_OP_94J1_122_9915_n209 DP_OP_94J1_122_9915_n205 DP_OP_94J1_122_9915_n199 DP_OP_94J1_122_9915_n127 DP_OP_94J1_122_9915_n128 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U99 VSS VDD  DP_OP_94J1_122_9915_n207 DP_OP_94J1_122_9915_n203 DP_OP_94J1_122_9915_n201 DP_OP_94J1_122_9915_n125 DP_OP_94J1_122_9915_n126 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U97 VSS VDD  DP_OP_94J1_122_9915_n189 DP_OP_94J1_122_9915_n195 DP_OP_94J1_122_9915_n122 DP_OP_94J1_122_9915_n123 DP_OP_94J1_122_9915_n124 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U95 VSS VDD  DP_OP_94J1_122_9915_n150 DP_OP_94J1_122_9915_n136 DP_OP_94J1_122_9915_n119 DP_OP_94J1_122_9915_n120 DP_OP_94J1_122_9915_n121 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U94 VSS VDD  DP_OP_94J1_122_9915_n148 DP_OP_94J1_122_9915_n142 DP_OP_94J1_122_9915_n146 DP_OP_94J1_122_9915_n117 DP_OP_94J1_122_9915_n118 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U93 VSS VDD  DP_OP_94J1_122_9915_n152 DP_OP_94J1_122_9915_n154 DP_OP_94J1_122_9915_n144 DP_OP_94J1_122_9915_n115 DP_OP_94J1_122_9915_n116 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U91 VSS VDD  DP_OP_94J1_122_9915_n192 DP_OP_94J1_122_9915_n134 DP_OP_94J1_122_9915_n112 DP_OP_94J1_122_9915_n113 DP_OP_94J1_122_9915_n114 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U89 VSS VDD  DP_OP_94J1_122_9915_n182 DP_OP_94J1_122_9915_n179 DP_OP_94J1_122_9915_n109 DP_OP_94J1_122_9915_n110 DP_OP_94J1_122_9915_n111 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U88 VSS VDD  DP_OP_94J1_122_9915_n128 DP_OP_94J1_122_9915_n177 DP_OP_94J1_122_9915_n131 DP_OP_94J1_122_9915_n107 DP_OP_94J1_122_9915_n108 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U86 VSS VDD  DP_OP_94J1_122_9915_n116 DP_OP_94J1_122_9915_n126 DP_OP_94J1_122_9915_n104 DP_OP_94J1_122_9915_n105 DP_OP_94J1_122_9915_n106 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U84 VSS VDD  DP_OP_94J1_122_9915_n170 DP_OP_94J1_122_9915_n124 DP_OP_94J1_122_9915_n101 DP_OP_94J1_122_9915_n102 DP_OP_94J1_122_9915_n103 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U82 VSS VDD  DP_OP_94J1_122_9915_n172 DP_OP_94J1_122_9915_n114 DP_OP_94J1_122_9915_n98 DP_OP_94J1_122_9915_n99 DP_OP_94J1_122_9915_n100 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U80 VSS VDD  DP_OP_94J1_122_9915_n111 DP_OP_94J1_122_9915_n108 DP_OP_94J1_122_9915_n95 DP_OP_94J1_122_9915_n96 DP_OP_94J1_122_9915_n97 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U78 VSS VDD  DP_OP_94J1_122_9915_n106 DP_OP_94J1_122_9915_n165 DP_OP_94J1_122_9915_n92 DP_OP_94J1_122_9915_n93 DP_OP_94J1_122_9915_n94 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U77 VSS VDD  DP_OP_94J1_122_9915_n100 DP_OP_94J1_122_9915_n103 DP_OP_94J1_122_9915_n160 DP_OP_94J1_122_9915_n90 DP_OP_94J1_122_9915_n91 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U75 VSS VDD  DP_OP_94J1_122_9915_n94 DP_OP_94J1_122_9915_n97 DP_OP_94J1_122_9915_n87 DP_OP_94J1_122_9915_n88 DP_OP_94J1_122_9915_n89 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U69 VSS VDD  DP_OP_94J1_122_9915_n151 DP_OP_94J1_122_9915_n137 DP_OP_94J1_122_9915_n149 DP_OP_94J1_122_9915_n80 DP_OP_94J1_122_9915_n81 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U68 VSS VDD  DP_OP_94J1_122_9915_n147 DP_OP_94J1_122_9915_n143 DP_OP_94J1_122_9915_n135 DP_OP_94J1_122_9915_n78 DP_OP_94J1_122_9915_n79 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U67 VSS VDD  DP_OP_94J1_122_9915_n139 DP_OP_94J1_122_9915_n141 DP_OP_94J1_122_9915_n145 DP_OP_94J1_122_9915_n76 DP_OP_94J1_122_9915_n77 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U66 VSS VDD  DP_OP_94J1_122_9915_n125 DP_OP_94J1_122_9915_n133 DP_OP_94J1_122_9915_n130 DP_OP_94J1_122_9915_n74 DP_OP_94J1_122_9915_n75 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U65 VSS VDD  DP_OP_94J1_122_9915_n84 DP_OP_94J1_122_9915_n127 DP_OP_94J1_122_9915_n115 DP_OP_94J1_122_9915_n72 DP_OP_94J1_122_9915_n73 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U63 VSS VDD  DP_OP_94J1_122_9915_n120 DP_OP_94J1_122_9915_n77 DP_OP_94J1_122_9915_n69 DP_OP_94J1_122_9915_n70 DP_OP_94J1_122_9915_n71 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U62 VSS VDD  DP_OP_94J1_122_9915_n81 DP_OP_94J1_122_9915_n117 DP_OP_94J1_122_9915_n79 DP_OP_94J1_122_9915_n67 DP_OP_94J1_122_9915_n68 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U61 VSS VDD  DP_OP_94J1_122_9915_n75 DP_OP_94J1_122_9915_n113 DP_OP_94J1_122_9915_n107 DP_OP_94J1_122_9915_n65 DP_OP_94J1_122_9915_n66 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U60 VSS VDD  DP_OP_94J1_122_9915_n73 DP_OP_94J1_122_9915_n110 DP_OP_94J1_122_9915_n105 DP_OP_94J1_122_9915_n63 DP_OP_94J1_122_9915_n64 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U58 VSS VDD  DP_OP_94J1_122_9915_n71 DP_OP_94J1_122_9915_n68 DP_OP_94J1_122_9915_n60 DP_OP_94J1_122_9915_n61 DP_OP_94J1_122_9915_n62 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U57 VSS VDD  DP_OP_94J1_122_9915_n66 DP_OP_94J1_122_9915_n99 DP_OP_94J1_122_9915_n96 DP_OP_94J1_122_9915_n58 DP_OP_94J1_122_9915_n59 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U56 VSS VDD  DP_OP_94J1_122_9915_n93 DP_OP_94J1_122_9915_n64 DP_OP_94J1_122_9915_n62 DP_OP_94J1_122_9915_n56 DP_OP_94J1_122_9915_n57 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U55 VSS VDD  DP_OP_94J1_122_9915_n59 DP_OP_94J1_122_9915_n90 DP_OP_94J1_122_9915_n88 DP_OP_94J1_122_9915_n54 DP_OP_94J1_122_9915_n55 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U53 VSS VDD  DP_OP_94J1_122_9915_n76 DP_OP_94J1_122_9915_n83 DP_OP_94J1_122_9915_n80 DP_OP_94J1_122_9915_n51 DP_OP_94J1_122_9915_n52 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U51 VSS VDD  DP_OP_94J1_122_9915_n74 DP_OP_94J1_122_9915_n72 DP_OP_94J1_122_9915_n48 DP_OP_94J1_122_9915_n49 DP_OP_94J1_122_9915_n50 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U50 VSS VDD  DP_OP_94J1_122_9915_n67 DP_OP_94J1_122_9915_n52 DP_OP_94J1_122_9915_n70 DP_OP_94J1_122_9915_n46 DP_OP_94J1_122_9915_n47 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U49 VSS VDD  DP_OP_94J1_122_9915_n50 DP_OP_94J1_122_9915_n65 DP_OP_94J1_122_9915_n63 DP_OP_94J1_122_9915_n44 DP_OP_94J1_122_9915_n45 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U47 VSS VDD  DP_OP_94J1_122_9915_n61 DP_OP_94J1_122_9915_n47 DP_OP_94J1_122_9915_n41 DP_OP_94J1_122_9915_n42 DP_OP_94J1_122_9915_n43 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U46 VSS VDD  DP_OP_94J1_122_9915_n56 DP_OP_94J1_122_9915_n45 DP_OP_94J1_122_9915_n43 DP_OP_94J1_122_9915_n39 DP_OP_94J1_122_9915_n40 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U44 VSS VDD  DP_OP_94J1_122_9915_n49 DP_OP_94J1_122_9915_n46 DP_OP_94J1_122_9915_n36 DP_OP_94J1_122_9915_n37 DP_OP_94J1_122_9915_n38 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U43 VSS VDD  DP_OP_94J1_122_9915_n38 DP_OP_94J1_122_9915_n44 DP_OP_94J1_122_9915_n42 DP_OP_94J1_122_9915_n34 DP_OP_94J1_122_9915_n35 FAx1_ASAP7_75t_R
XU3 VSS VDD  n14 n6 INVx2_ASAP7_75t_R
XU4 VSS VDD  DP_OP_94J1_122_9915_n153 n26 DP_OP_94J1_122_9915_n84 XOR2xp5_ASAP7_75t_R
XU5 VSS VDD  n5 TIEHIx1_ASAP7_75t_R
XU6 VSS VDD  n5 out[9] INVx1_ASAP7_75t_R
XU7 VSS VDD  n5 out[10] INVx1_ASAP7_75t_R
XU8 VSS VDD  n5 out[11] INVx1_ASAP7_75t_R
XU9 VSS VDD  n5 out[12] INVx1_ASAP7_75t_R
XU10 VSS VDD  n8 n17 INVx3_ASAP7_75t_R
XU11 VSS VDD  DP_OP_94J1_122_9915_n159 n14 BUFx4_ASAP7_75t_R
XU12 VSS VDD  DP_OP_94J1_122_9915_n222 n8 BUFx4_ASAP7_75t_R
XU13 VSS VDD  DP_OP_94J1_122_9915_n55 n7 BUFx4_ASAP7_75t_R
XU14 VSS VDD  n7 n13 INVx4_ASAP7_75t_R
XU15 VSS VDD  in[7] in[15] n26 NAND2xp33_ASAP7_75t_R
XU16 VSS VDD  DP_OP_94J1_122_9915_n153 n26 DP_OP_94J1_122_9915_n83 NOR2x1_ASAP7_75t_R
XU17 VSS VDD  in[12] in[20] DP_OP_94J1_122_9915_n246 NAND2xp5_ASAP7_75t_R
XU18 VSS VDD  in[5] in[13] DP_OP_94J1_122_9915_n194 NAND2xp5_ASAP7_75t_R
XU19 VSS VDD  in[6] in[14] DP_OP_94J1_122_9915_n132 NAND2xp5_ASAP7_75t_R
XU20 VSS VDD  DP_OP_94J1_122_9915_n34 n25 INVxp67_ASAP7_75t_R
XU21 VSS VDD  n11 DP_OP_94J1_122_9915_n40 DP_OP_94J1_122_9915_n54 n9 MAJIxp5_ASAP7_75t_R
XU22 VSS VDD  n12 DP_OP_94J1_122_9915_n39 DP_OP_94J1_122_9915_n35 n10 MAJIxp5_ASAP7_75t_R
XU23 VSS VDD  n13 n22 DP_OP_94J1_122_9915_n57 n11 MAJIxp5_ASAP7_75t_R
XU24 VSS VDD  n13 n22 DP_OP_94J1_122_9915_n57 n23 MAJx2_ASAP7_75t_R
XU25 VSS VDD  n12 DP_OP_94J1_122_9915_n39 DP_OP_94J1_122_9915_n35 n24 MAJx2_ASAP7_75t_R
XU26 VSS VDD  n11 DP_OP_94J1_122_9915_n40 DP_OP_94J1_122_9915_n54 n12 MAJx2_ASAP7_75t_R
XU27 VSS VDD  DP_OP_94J1_122_9915_n292 DP_OP_94J1_122_9915_n294 DP_OP_94J1_122_9915_n296 A0  n15 FAx1_ASAP7_75t_R
XU28 VSS VDD  DP_OP_94J1_122_9915_n275 n16 INVx1_ASAP7_75t_R
XU29 VSS VDD  DP_OP_94J1_122_9915_n38 DP_OP_94J1_122_9915_n44 DP_OP_94J1_122_9915_n42 n18 MAJIxp5_ASAP7_75t_R
XU30 VSS VDD  DP_OP_94J1_122_9915_n158 DP_OP_94J1_122_9915_n87 INVx1_ASAP7_75t_R
XU31 VSS VDD  DP_OP_94J1_122_9915_n272 DP_OP_94J1_122_9915_n220 INVx1_ASAP7_75t_R
XU32 VSS VDD  DP_OP_94J1_122_9915_n280 DP_OP_94J1_122_9915_n271 INVx1_ASAP7_75t_R
XU33 VSS VDD  DP_OP_94J1_122_9915_n232 DP_OP_94J1_122_9915_n223 INVx1_ASAP7_75t_R
XU34 VSS VDD  DP_OP_94J1_122_9915_n162 DP_OP_94J1_122_9915_n92 INVx1_ASAP7_75t_R
XU35 VSS VDD  DP_OP_94J1_122_9915_n186 DP_OP_94J1_122_9915_n164 INVx1_ASAP7_75t_R
XU36 VSS VDD  DP_OP_94J1_122_9915_n58 DP_OP_94J1_122_9915_n41 INVx1_ASAP7_75t_R
XU37 VSS VDD  DP_OP_94J1_122_9915_n168 DP_OP_94J1_122_9915_n95 INVx1_ASAP7_75t_R
XU38 VSS VDD  DP_OP_94J1_122_9915_n268 DP_OP_94J1_122_9915_n230 INVx1_ASAP7_75t_R
XU39 VSS VDD  DP_OP_94J1_122_9915_n183 DP_OP_94J1_122_9915_n167 INVx1_ASAP7_75t_R
XU40 VSS VDD  DP_OP_94J1_122_9915_n121 DP_OP_94J1_122_9915_n98 INVx1_ASAP7_75t_R
XU41 VSS VDD  DP_OP_94J1_122_9915_n102 DP_OP_94J1_122_9915_n60 INVx1_ASAP7_75t_R
XU42 VSS VDD  DP_OP_94J1_122_9915_n118 DP_OP_94J1_122_9915_n101 INVx1_ASAP7_75t_R
XU43 VSS VDD  DP_OP_94J1_122_9915_n175 DP_OP_94J1_122_9915_n104 INVx1_ASAP7_75t_R
XU44 VSS VDD  DP_OP_94J1_122_9915_n208 DP_OP_94J1_122_9915_n174 INVx1_ASAP7_75t_R
XU45 VSS VDD  DP_OP_94J1_122_9915_n185 DP_OP_94J1_122_9915_n109 INVx1_ASAP7_75t_R
XU46 VSS VDD  DP_OP_94J1_122_9915_n198 DP_OP_94J1_122_9915_n184 INVx1_ASAP7_75t_R
XU47 VSS VDD  DP_OP_94J1_122_9915_n239 DP_OP_94J1_122_9915_n181 INVx1_ASAP7_75t_R
XU48 VSS VDD  DP_OP_94J1_122_9915_n138 DP_OP_94J1_122_9915_n112 INVx1_ASAP7_75t_R
XU49 VSS VDD  DP_OP_94J1_122_9915_n123 DP_OP_94J1_122_9915_n69 INVx1_ASAP7_75t_R
XU50 VSS VDD  DP_OP_94J1_122_9915_n140 DP_OP_94J1_122_9915_n122 INVx1_ASAP7_75t_R
XU51 VSS VDD  DP_OP_94J1_122_9915_n187 DP_OP_94J1_122_9915_n119 INVx1_ASAP7_75t_R
XU52 VSS VDD  DP_OP_94J1_122_9915_n51 DP_OP_94J1_122_9915_n36 INVx1_ASAP7_75t_R
XU53 VSS VDD  DP_OP_94J1_122_9915_n78 DP_OP_94J1_122_9915_n48 INVx1_ASAP7_75t_R
XU54 VSS VDD  in[7] in[15] A1  DP_OP_94J1_122_9915_n129 HAxp5_ASAP7_75t_R
XU55 VSS VDD  in[6] in[14] A2  DP_OP_94J1_122_9915_n191 HAxp5_ASAP7_75t_R
XU56 VSS VDD  in[5] in[13] A3  DP_OP_94J1_122_9915_n243 HAxp5_ASAP7_75t_R
XU57 VSS VDD  in[12] in[20] A4  DP_OP_94J1_122_9915_n278 HAxp5_ASAP7_75t_R
XU58 VSS VDD  DP_OP_94J1_122_9915_n273 DP_OP_94J1_122_9915_n277 n16 A5  out[0] FAx1_ASAP7_75t_R
XU59 VSS VDD  n15 DP_OP_94J1_122_9915_n277 DP_OP_94J1_122_9915_n273 n19 MAJIxp5_ASAP7_75t_R
XU60 VSS VDD  DP_OP_94J1_122_9915_n225 n19 n17 A6  out[1] FAx1_ASAP7_75t_R
XU61 VSS VDD  n17 n19 DP_OP_94J1_122_9915_n225 n20 MAJIxp5_ASAP7_75t_R
XU62 VSS VDD  DP_OP_94J1_122_9915_n161 n20 n14 A7  out[2] FAx1_ASAP7_75t_R
XU63 VSS VDD  n6 n20 DP_OP_94J1_122_9915_n161 n21 MAJIxp5_ASAP7_75t_R
XU64 VSS VDD  DP_OP_94J1_122_9915_n91 DP_OP_94J1_122_9915_n89 n21 A8  out[3] FAx1_ASAP7_75t_R
XU65 VSS VDD  DP_OP_94J1_122_9915_n91 DP_OP_94J1_122_9915_n89 n21 n22 MAJx2_ASAP7_75t_R
XU66 VSS VDD  DP_OP_94J1_122_9915_n57 n22 n13 A9  out[4] FAx1_ASAP7_75t_R
XU67 VSS VDD  DP_OP_94J1_122_9915_n54 DP_OP_94J1_122_9915_n40 n23 A10  out[5] FAx1_ASAP7_75t_R
XU68 VSS VDD  DP_OP_94J1_122_9915_n35 DP_OP_94J1_122_9915_n39 n9 A11  out[6] FAx1_ASAP7_75t_R
XU69 VSS VDD  n18 DP_OP_94J1_122_9915_n37 n24 A12  out[7] FAx1_ASAP7_75t_R
XU70 VSS VDD  n25 DP_OP_94J1_122_9915_n37 n10 out[8] MAJIxp5_ASAP7_75t_R
.ENDS


