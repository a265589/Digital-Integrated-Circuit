.SUBCKT Control VSS VDD  clk rst_n out_valid
Xcounter_reg_0_ VSS VDD clk N_8  n4 n13 n7 ASYNC_DFFHx1_ASAP7_75t_R
Xcounter_reg_2_ VSS VDD clk  N_10 n4 n8 n6 ASYNC_DFFHx1_ASAP7_75t_R
Xcounter_reg_1_ VSS VDD clk  N_9 n4 n12 n5 ASYNC_DFFHx1_ASAP7_75t_R
Xout_valid_reg VSS VDD  clk N_12 n4 n11 n3 ASYNC_DFFHx1_ASAP7_75t_R
XU12 VSS VDD  n6 n10 BUFx5_ASAP7_75t_R
XU13 VSS VDD  n7 n5 n9 NAND2xp33_ASAP7_75t_R
XU14 VSS VDD  n7 n5 n14 AND2x2_ASAP7_75t_R
XU15 VSS VDD  n10 n16 INVx2_ASAP7_75t_R
XU16 VSS VDD  rst_n n11 INVx8_ASAP7_75t_R
XU17 VSS VDD  rst_n n12 INVx8_ASAP7_75t_R
XU18 VSS VDD  rst_n n13 INVx8_ASAP7_75t_R
XU19 VSS VDD  rst_n n8 INVx8_ASAP7_75t_R
XU20 VSS VDD  n4 TIELOx1_ASAP7_75t_R
XU21 VSS VDD  n3 out_valid INVxp33_ASAP7_75t_R
XU22 VSS VDD  n10 n9 N_12 NOR2xp33_ASAP7_75t_R
XU23 VSS VDD  n7 n5 n15 NOR2xp33_ASAP7_75t_R
XU24 VSS VDD  n15 n16 n14 N_9 NOR3xp33_ASAP7_75t_R
XU25 VSS VDD  n10 n7 N_8 AND2x2_ASAP7_75t_R
XU26 VSS VDD  n7 n16 n5 N_10 NOR3xp33_ASAP7_75t_R
.ENDS


