.SUBCKT Accumulator VSS VDD  clk rst_n in_valid partial_sum[12] partial_sum[11] partial_sum[10] partial_sum[9] partial_sum[8] partial_sum[7] partial_sum[6] partial_sum[5] partial_sum[4] partial_sum[3] partial_sum[2] partial_sum[1] partial_sum[0] result[12] result[11] result[10] result[9] result[8] result[7] result[6] result[5] result[4] result[3] result[2] result[1] result[0]
Xresult_reg_12_ VSS VDD  n54 clk n29 n98 n53 ASYNC_DFFHx1_ASAP7_75t_R
Xresult_reg_11_ VSS VDD  n52 clk n29 n96 n51 ASYNC_DFFHx1_ASAP7_75t_R
Xresult_reg_10_ VSS VDD  n50 clk n29 n69 n49 ASYNC_DFFHx1_ASAP7_75t_R
Xresult_reg_9_ VSS VDD  n48 clk n29 n64 n47 ASYNC_DFFHx1_ASAP7_75t_R
Xresult_reg_8_ VSS VDD  n46 clk n29 n72 n45 ASYNC_DFFHx1_ASAP7_75t_R
Xresult_reg_7_ VSS VDD  n44 clk n29 n67 n43 ASYNC_DFFHx1_ASAP7_75t_R
Xresult_reg_6_ VSS VDD  n42 clk n29 n66 n41 ASYNC_DFFHx1_ASAP7_75t_R
Xresult_reg_5_ VSS VDD  n40 clk n29 n68 n39 ASYNC_DFFHx1_ASAP7_75t_R
Xresult_reg_4_ VSS VDD  n38 clk n29 n97 n37 ASYNC_DFFHx1_ASAP7_75t_R
Xresult_reg_3_ VSS VDD  n36 clk n29 n55 n35 ASYNC_DFFHx1_ASAP7_75t_R
Xresult_reg_2_ VSS VDD  n34 clk n29 n65 n33 ASYNC_DFFHx1_ASAP7_75t_R
Xresult_reg_1_ VSS VDD  n32 clk n29 n71 n31 ASYNC_DFFHx1_ASAP7_75t_R
Xresult_reg_0_ VSS VDD  n30 clk n29 n95 n28 ASYNC_DFFHx1_ASAP7_75t_R
XU57 VSS VDD  n182 result[12] INVx1_ASAP7_75t_R
XU58 VSS VDD  n82 result[1] INVx1_ASAP7_75t_R
XU59 VSS VDD  n189 result[0] INVx3_ASAP7_75t_R
XU60 VSS VDD  n188 result[2] INVx4_ASAP7_75t_R
XU61 VSS VDD  n185 result[8] INVx4_ASAP7_75t_R
XU62 VSS VDD  n184 result[10] INVx4_ASAP7_75t_R
XU63 VSS VDD  n186 result[6] INVx4_ASAP7_75t_R
XU64 VSS VDD  n187 result[4] INVx4_ASAP7_75t_R
XU65 VSS VDD  n35 n74 BUFx5_ASAP7_75t_R
XU66 VSS VDD  n39 n75 BUFx5_ASAP7_75t_R
XU67 VSS VDD  n43 n76 BUFx5_ASAP7_75t_R
XU68 VSS VDD  n47 n77 BUFx5_ASAP7_75t_R
XU69 VSS VDD  in_valid n56 INVx8_ASAP7_75t_R
XU70 VSS VDD  in_valid n57 INVx8_ASAP7_75t_R
XU71 VSS VDD  in_valid n58 INVx8_ASAP7_75t_R
XU72 VSS VDD  in_valid n59 INVx8_ASAP7_75t_R
XU73 VSS VDD  in_valid n60 INVx8_ASAP7_75t_R
XU74 VSS VDD  in_valid n61 INVx8_ASAP7_75t_R
XU75 VSS VDD  in_valid n62 INVx8_ASAP7_75t_R
XU76 VSS VDD  in_valid n63 INVx8_ASAP7_75t_R
XU77 VSS VDD  rst_n n64 INVx8_ASAP7_75t_R
XU78 VSS VDD  rst_n n65 INVx8_ASAP7_75t_R
XU79 VSS VDD  rst_n n66 INVx8_ASAP7_75t_R
XU80 VSS VDD  rst_n n67 INVx8_ASAP7_75t_R
XU81 VSS VDD  rst_n n68 INVx8_ASAP7_75t_R
XU82 VSS VDD  rst_n n69 INVx8_ASAP7_75t_R
XU83 VSS VDD  n31 n82 BUFx5_ASAP7_75t_R
XU84 VSS VDD  rst_n n71 INVx8_ASAP7_75t_R
XU85 VSS VDD  rst_n n72 INVx8_ASAP7_75t_R
XU86 VSS VDD  n53 n182 BUFx5_ASAP7_75t_R
XU87 VSS VDD  n74 result[3] INVx2_ASAP7_75t_R
XU88 VSS VDD  n75 result[5] INVx2_ASAP7_75t_R
XU89 VSS VDD  n76 result[7] INVx2_ASAP7_75t_R
XU90 VSS VDD  n77 result[9] INVx2_ASAP7_75t_R
XU91 VSS VDD  n49 n184 BUFx5_ASAP7_75t_R
XU92 VSS VDD  n51 n183 BUFx5_ASAP7_75t_R
XU93 VSS VDD  n183 result[11] INVx4_ASAP7_75t_R
XU94 VSS VDD  n28 n189 BUFx5_ASAP7_75t_R
XU95 VSS VDD  n41 n186 BUFx5_ASAP7_75t_R
XU96 VSS VDD  n37 n187 BUFx5_ASAP7_75t_R
XU97 VSS VDD  n33 n188 BUFx5_ASAP7_75t_R
XU98 VSS VDD  n45 n185 BUFx5_ASAP7_75t_R
XU99 VSS VDD  partial_sum[2] n99 INVx8_ASAP7_75t_R
XU100 VSS VDD  partial_sum[10] n87 INVx8_ASAP7_75t_R
XU101 VSS VDD  partial_sum[10] n162 INVx8_ASAP7_75t_R
XU102 VSS VDD  partial_sum[8] n88 INVx8_ASAP7_75t_R
XU103 VSS VDD  partial_sum[8] n121 INVx8_ASAP7_75t_R
XU104 VSS VDD  partial_sum[6] n89 INVx8_ASAP7_75t_R
XU105 VSS VDD  partial_sum[6] n154 INVx8_ASAP7_75t_R
XU106 VSS VDD  partial_sum[4] n90 INVx8_ASAP7_75t_R
XU107 VSS VDD  partial_sum[4] n106 INVx8_ASAP7_75t_R
XU108 VSS VDD  in_valid n91 INVx8_ASAP7_75t_R
XU109 VSS VDD  in_valid n92 INVx8_ASAP7_75t_R
XU110 VSS VDD  in_valid n93 INVx8_ASAP7_75t_R
XU111 VSS VDD  in_valid n94 INVx8_ASAP7_75t_R
XU112 VSS VDD  in_valid n179 INVx8_ASAP7_75t_R
XU113 VSS VDD  rst_n n95 INVx8_ASAP7_75t_R
XU114 VSS VDD  rst_n n96 INVx8_ASAP7_75t_R
XU115 VSS VDD  rst_n n97 INVx8_ASAP7_75t_R
XU116 VSS VDD  rst_n n98 INVx8_ASAP7_75t_R
XU117 VSS VDD  rst_n n55 INVx8_ASAP7_75t_R
XU118 VSS VDD  n29 TIELOx1_ASAP7_75t_R
XU119 VSS VDD  result[0] partial_sum[1] n170 NAND2xp33_ASAP7_75t_R
XU120 VSS VDD  n99 n170 n82 n132 MAJIxp5_ASAP7_75t_R
XU121 VSS VDD  result[2] partial_sum[3] n132 n110 MAJIxp5_ASAP7_75t_R
XU122 VSS VDD  n74 n110 n90 n117 MAJIxp5_ASAP7_75t_R
XU123 VSS VDD  result[4] partial_sum[5] n117 n158 MAJIxp5_ASAP7_75t_R
XU124 VSS VDD  n75 n158 n89 n139 MAJIxp5_ASAP7_75t_R
XU125 VSS VDD  result[6] partial_sum[7] n139 n122 MAJIxp5_ASAP7_75t_R
XU126 VSS VDD  n76 n121 n101 NOR2xp33_ASAP7_75t_R
XU127 VSS VDD  result[7] partial_sum[8] n100 NOR2xp33_ASAP7_75t_R
XU128 VSS VDD  n101 n100 n102 NOR2xp33_ASAP7_75t_R
XU129 VSS VDD  n122 n102 A0  n103 HAxp5_ASAP7_75t_R
XU130 VSS VDD  in_valid n103 n105 NAND2xp33_ASAP7_75t_R
XU131 VSS VDD  result[8] n57 n104 NAND2xp33_ASAP7_75t_R
XU132 VSS VDD  n105 n104 n46 NAND2xp33_ASAP7_75t_R
XU133 VSS VDD  n74 n106 n108 NOR2xp33_ASAP7_75t_R
XU134 VSS VDD  result[3] partial_sum[4] n107 NOR2xp33_ASAP7_75t_R
XU135 VSS VDD  n108 n107 n109 NOR2xp33_ASAP7_75t_R
XU136 VSS VDD  n110 n109 A1  n111 HAxp5_ASAP7_75t_R
XU137 VSS VDD  in_valid n111 n113 NAND2xp33_ASAP7_75t_R
XU138 VSS VDD  result[4] n58 n112 NAND2xp33_ASAP7_75t_R
XU139 VSS VDD  n113 n112 n38 NAND2xp33_ASAP7_75t_R
XU140 VSS VDD  result[4] partial_sum[5] n115 NAND2xp33_ASAP7_75t_R
XU141 VSS VDD  result[4] partial_sum[5] n114 OR2x2_ASAP7_75t_R
XU142 VSS VDD  n115 n114 n116 NAND2xp33_ASAP7_75t_R
XU143 VSS VDD  n117 n116 A2  n118 HAxp5_ASAP7_75t_R
XU144 VSS VDD  in_valid n118 n120 NAND2xp33_ASAP7_75t_R
XU145 VSS VDD  result[5] n60 n119 NAND2xp33_ASAP7_75t_R
XU146 VSS VDD  n120 n119 n40 NAND2xp33_ASAP7_75t_R
XU147 VSS VDD  n76 n122 n88 n143 MAJIxp5_ASAP7_75t_R
XU148 VSS VDD  result[8] partial_sum[9] n124 NAND2xp33_ASAP7_75t_R
XU149 VSS VDD  result[8] partial_sum[9] n123 OR2x2_ASAP7_75t_R
XU150 VSS VDD  n124 n123 n125 NAND2xp33_ASAP7_75t_R
XU151 VSS VDD  n143 n125 A3  n126 HAxp5_ASAP7_75t_R
XU152 VSS VDD  in_valid n126 n128 NAND2xp33_ASAP7_75t_R
XU153 VSS VDD  result[9] n61 n127 NAND2xp33_ASAP7_75t_R
XU154 VSS VDD  n128 n127 n48 NAND2xp33_ASAP7_75t_R
XU155 VSS VDD  result[2] partial_sum[3] n130 NAND2xp33_ASAP7_75t_R
XU156 VSS VDD  result[2] partial_sum[3] n129 OR2x2_ASAP7_75t_R
XU157 VSS VDD  n130 n129 n131 NAND2xp33_ASAP7_75t_R
XU158 VSS VDD  n132 n131 A4  n133 HAxp5_ASAP7_75t_R
XU159 VSS VDD  in_valid n133 n135 NAND2xp33_ASAP7_75t_R
XU160 VSS VDD  result[3] n56 n134 NAND2xp33_ASAP7_75t_R
XU161 VSS VDD  n135 n134 n36 NAND2xp33_ASAP7_75t_R
XU162 VSS VDD  result[6] partial_sum[7] n137 NAND2xp33_ASAP7_75t_R
XU163 VSS VDD  result[6] partial_sum[7] n136 OR2x2_ASAP7_75t_R
XU164 VSS VDD  n137 n136 n138 NAND2xp33_ASAP7_75t_R
XU165 VSS VDD  n139 n138 A5  n140 HAxp5_ASAP7_75t_R
XU166 VSS VDD  in_valid n140 n142 NAND2xp33_ASAP7_75t_R
XU167 VSS VDD  result[7] n62 n141 NAND2xp33_ASAP7_75t_R
XU168 VSS VDD  n142 n141 n44 NAND2xp33_ASAP7_75t_R
XU169 VSS VDD  result[8] partial_sum[9] n143 n163 MAJIxp5_ASAP7_75t_R
XU170 VSS VDD  n77 n162 n145 NOR2xp33_ASAP7_75t_R
XU171 VSS VDD  result[9] partial_sum[10] n144 NOR2xp33_ASAP7_75t_R
XU172 VSS VDD  n145 n144 n146 NOR2xp33_ASAP7_75t_R
XU173 VSS VDD  n163 n146 A6  n147 HAxp5_ASAP7_75t_R
XU174 VSS VDD  in_valid n147 n149 NAND2xp33_ASAP7_75t_R
XU175 VSS VDD  result[10] n92 n148 NAND2xp33_ASAP7_75t_R
XU176 VSS VDD  n149 n148 n50 NAND2xp33_ASAP7_75t_R
XU177 VSS VDD  partial_sum[2] n170 A7  n150 HAxp5_ASAP7_75t_R
XU178 VSS VDD  n150 n82 A8  n151 HAxp5_ASAP7_75t_R
XU179 VSS VDD  in_valid n151 n153 NAND2xp33_ASAP7_75t_R
XU180 VSS VDD  result[2] n59 n152 NAND2xp33_ASAP7_75t_R
XU181 VSS VDD  n153 n152 n34 NAND2xp33_ASAP7_75t_R
XU182 VSS VDD  n75 n154 n156 NOR2xp33_ASAP7_75t_R
XU183 VSS VDD  result[5] partial_sum[6] n155 NOR2xp33_ASAP7_75t_R
XU184 VSS VDD  n156 n155 n157 NOR2xp33_ASAP7_75t_R
XU185 VSS VDD  n158 n157 A9  n159 HAxp5_ASAP7_75t_R
XU186 VSS VDD  in_valid n159 n161 NAND2xp33_ASAP7_75t_R
XU187 VSS VDD  result[6] n63 n160 NAND2xp33_ASAP7_75t_R
XU188 VSS VDD  n161 n160 n42 NAND2xp33_ASAP7_75t_R
XU189 VSS VDD  n77 n163 n87 n176 MAJIxp5_ASAP7_75t_R
XU190 VSS VDD  result[10] partial_sum[11] n165 OR2x2_ASAP7_75t_R
XU191 VSS VDD  result[10] partial_sum[11] n164 NAND2xp33_ASAP7_75t_R
XU192 VSS VDD  n165 n164 n166 NAND2xp33_ASAP7_75t_R
XU193 VSS VDD  n176 n166 A10  n167 HAxp5_ASAP7_75t_R
XU194 VSS VDD  in_valid n167 n169 NAND2xp33_ASAP7_75t_R
XU195 VSS VDD  result[11] n179 n168 NAND2xp33_ASAP7_75t_R
XU196 VSS VDD  n169 n168 n52 NAND2xp33_ASAP7_75t_R
XU197 VSS VDD  result[0] partial_sum[1] n171 OR2x2_ASAP7_75t_R
XU198 VSS VDD  n171 in_valid n170 n173 NAND3xp33_ASAP7_75t_R
XU199 VSS VDD  result[1] n93 n172 NAND2xp33_ASAP7_75t_R
XU200 VSS VDD  n173 n172 n32 NAND2xp33_ASAP7_75t_R
XU201 VSS VDD  in_valid partial_sum[0] n175 NAND2xp33_ASAP7_75t_R
XU202 VSS VDD  result[0] n91 n174 NAND2xp33_ASAP7_75t_R
XU203 VSS VDD  n175 n174 n30 NAND2xp33_ASAP7_75t_R
XU204 VSS VDD  result[10] partial_sum[11] n176 n177 MAJIxp5_ASAP7_75t_R
XU205 VSS VDD  partial_sum[12] n177 result[11] A11  n178 FAx1_ASAP7_75t_R
XU206 VSS VDD  in_valid n178 n181 NAND2xp33_ASAP7_75t_R
XU207 VSS VDD  result[12] n94 n180 NAND2xp33_ASAP7_75t_R
XU208 VSS VDD  n181 n180 n54 NAND2xp33_ASAP7_75t_R
.ENDS


