.TITLE DIC_Final

***-----------------------***
***        setting        ***
***-----------------------***

.protect
.include '../08_TECH/LIB/7nm_TT.pm'
.include '../08_TECH/LIB/16mos.pm'
.include '../08_TECH/LIB/asap7sc7p5t_SIMPLE_RVT.sp' 
.include '../08_TECH/LIB/asap7sc7p5t_SEQ_RVT.sp'    
.include '../08_TECH/LIB/asap7sc7p5t_INVBUF_RVT.sp' 
.include '../08_TECH/LIB/asap7sc7p5t_AO_RVT.sp'     
.include '../08_TECH/LIB/asap7sc7p5t_OA_RVT.sp'     
.unprotect

.VEC "mul.vec" 

*** Voltage: 0.7V ***
.PARAM supply=0.7v

*** Temperature: 25C ***
.TEMP 25

***********************************
* Transition Analysis             *
***********************************
.TRAN 1ps 20ns 

***********************************
* HSPICE Options                  *
***********************************
.OPTION POST PROBE
.OPTION NOMOD BRIEF MEASDGT=7 
.OPTION CAPTAB NOTOP AUTOSTOP

***********************************
* Output Signals                  *
***********************************
.probe tran v(*) i(*)


***********************************
* Define Global Nets              *
***********************************
.GLOBAL VDD GND BL BLB

***********************************
* Voltage Sources                 *
***********************************
vdd     VDD   0  DC supply
vss     VSS   0  DC 0
vbl     BL    0   DC supply/2
vblb    BLB   0   DC supply/2

***********************************
* Measurement Commands            *
***********************************
.meas pwr avg POWER



***-----------------------***
***        circuit        ***
***-----------------------***


* // Xbuf Input In_bar INV
* // ADD INPUT BUFFER
* // WEIGHT IS INITIALIZE IN THE SRAM
* // SO CIM OPERATION IS READ THE WEIGHT AND THEN DO DOT PRODUCT 

X11 I111 O_1_1_1_1 WL_1_1 BL BLB W_1_1_1 W_1_1_1_bar CIM_cell
X12 I111 O_1_1_1_2 WL_1_1 BL BLB W_1_1_2 W_1_1_2_bar CIM_cell
X13 I111 O_1_1_1_3 WL_1_1 BL BLB W_1_1_3 W_1_1_3_bar CIM_cell
X14 I111 O_1_1_1_4 WL_1_1 BL BLB W_1_1_4 W_1_1_4_bar CIM_cell
X21 I112 O_1_1_2_1 WL_1_2 BL BLB W_1_1_1 W_1_1_1_bar CIM_cell
X22 I112 O_1_1_2_2 WL_1_2 BL BLB W_1_1_2 W_1_1_2_bar CIM_cell
X23 I112 O_1_1_2_3 WL_1_2 BL BLB W_1_1_3 W_1_1_3_bar CIM_cell
X24 I112 O_1_1_2_4 WL_1_2 BL BLB W_1_1_4 W_1_1_4_bar CIM_cell
X31 I113 O_1_1_3_1 WL_1_3 BL BLB W_1_1_1 W_1_1_1_bar CIM_cell
X32 I113 O_1_1_3_2 WL_1_3 BL BLB W_1_1_2 W_1_1_2_bar CIM_cell
X33 I113 O_1_1_3_3 WL_1_3 BL BLB W_1_1_3 W_1_1_3_bar CIM_cell
X34 I113 O_1_1_3_4 WL_1_3 BL BLB W_1_1_4 W_1_1_4_bar CIM_cell
X41 I114 O_1_1_4_1 WL_1_4 BL BLB W_1_1_1 W_1_1_1_bar CIM_cell
X42 I114 O_1_1_4_2 WL_1_4 BL BLB W_1_1_2 W_1_1_2_bar CIM_cell
X43 I114 O_1_1_4_3 WL_1_4 BL BLB W_1_1_3 W_1_1_3_bar CIM_cell
X44 I114 O_1_1_4_4 WL_1_4 BL BLB W_1_1_4 W_1_1_4_bar CIM_cell
X51 I121 O_1_2_1_1 WL_1_1 BL BLB W_1_2_1 W_1_2_1_bar CIM_cell
X52 I121 O_1_2_1_2 WL_1_1 BL BLB W_1_2_2 W_1_2_2_bar CIM_cell
X53 I121 O_1_2_1_3 WL_1_1 BL BLB W_1_2_3 W_1_2_3_bar CIM_cell
X54 I121 O_1_2_1_4 WL_1_1 BL BLB W_1_2_4 W_1_2_4_bar CIM_cell
X61 I122 O_1_2_2_1 WL_1_2 BL BLB W_1_2_1 W_1_2_1_bar CIM_cell
X62 I122 O_1_2_2_2 WL_1_2 BL BLB W_1_2_2 W_1_2_2_bar CIM_cell
X63 I122 O_1_2_2_3 WL_1_2 BL BLB W_1_2_3 W_1_2_3_bar CIM_cell
X64 I122 O_1_2_2_4 WL_1_2 BL BLB W_1_2_4 W_1_2_4_bar CIM_cell
X71 I123 O_1_2_3_1 WL_1_3 BL BLB W_1_2_1 W_1_2_1_bar CIM_cell
X72 I123 O_1_2_3_2 WL_1_3 BL BLB W_1_2_2 W_1_2_2_bar CIM_cell
X73 I123 O_1_2_3_3 WL_1_3 BL BLB W_1_2_3 W_1_2_3_bar CIM_cell
X74 I123 O_1_2_3_4 WL_1_3 BL BLB W_1_2_4 W_1_2_4_bar CIM_cell
X81 I124 O_1_2_4_1 WL_1_4 BL BLB W_1_2_1 W_1_2_1_bar CIM_cell
X82 I124 O_1_2_4_2 WL_1_4 BL BLB W_1_2_2 W_1_2_2_bar CIM_cell
X83 I124 O_1_2_4_3 WL_1_4 BL BLB W_1_2_3 W_1_2_3_bar CIM_cell
X84 I124 O_1_2_4_4 WL_1_4 BL BLB W_1_2_4 W_1_2_4_bar CIM_cell
X91 I131 O_1_3_1_1 WL_1_1 BL BLB W_1_3_1 W_1_3_1_bar CIM_cell
X92 I131 O_1_3_1_2 WL_1_1 BL BLB W_1_3_2 W_1_3_2_bar CIM_cell
X93 I131 O_1_3_1_3 WL_1_1 BL BLB W_1_3_3 W_1_3_3_bar CIM_cell
X94 I131 O_1_3_1_4 WL_1_1 BL BLB W_1_3_4 W_1_3_4_bar CIM_cell
X101 I132 O_1_3_2_1 WL_1_2 BL BLB W_1_3_1 W_1_3_1_bar CIM_cell
X102 I132 O_1_3_2_2 WL_1_2 BL BLB W_1_3_2 W_1_3_2_bar CIM_cell
X103 I132 O_1_3_2_3 WL_1_2 BL BLB W_1_3_3 W_1_3_3_bar CIM_cell
X104 I132 O_1_3_2_4 WL_1_2 BL BLB W_1_3_4 W_1_3_4_bar CIM_cell
X111 I133 O_1_3_3_1 WL_1_3 BL BLB W_1_3_1 W_1_3_1_bar CIM_cell
X112 I133 O_1_3_3_2 WL_1_3 BL BLB W_1_3_2 W_1_3_2_bar CIM_cell
X113 I133 O_1_3_3_3 WL_1_3 BL BLB W_1_3_3 W_1_3_3_bar CIM_cell
X114 I133 O_1_3_3_4 WL_1_3 BL BLB W_1_3_4 W_1_3_4_bar CIM_cell
X121 I134 O_1_3_4_1 WL_1_4 BL BLB W_1_3_1 W_1_3_1_bar CIM_cell
X122 I134 O_1_3_4_2 WL_1_4 BL BLB W_1_3_2 W_1_3_2_bar CIM_cell
X123 I134 O_1_3_4_3 WL_1_4 BL BLB W_1_3_3 W_1_3_3_bar CIM_cell
X124 I134 O_1_3_4_4 WL_1_4 BL BLB W_1_3_4 W_1_3_4_bar CIM_cell
X131 I141 O_1_4_1_1 WL_1_1 BL BLB W_1_4_1 W_1_4_1_bar CIM_cell
X132 I141 O_1_4_1_2 WL_1_1 BL BLB W_1_4_2 W_1_4_2_bar CIM_cell
X133 I141 O_1_4_1_3 WL_1_1 BL BLB W_1_4_3 W_1_4_3_bar CIM_cell
X134 I141 O_1_4_1_4 WL_1_1 BL BLB W_1_4_4 W_1_4_4_bar CIM_cell
X141 I142 O_1_4_2_1 WL_1_2 BL BLB W_1_4_1 W_1_4_1_bar CIM_cell
X142 I142 O_1_4_2_2 WL_1_2 BL BLB W_1_4_2 W_1_4_2_bar CIM_cell
X143 I142 O_1_4_2_3 WL_1_2 BL BLB W_1_4_3 W_1_4_3_bar CIM_cell
X144 I142 O_1_4_2_4 WL_1_2 BL BLB W_1_4_4 W_1_4_4_bar CIM_cell
X151 I143 O_1_4_3_1 WL_1_3 BL BLB W_1_4_1 W_1_4_1_bar CIM_cell
X152 I143 O_1_4_3_2 WL_1_3 BL BLB W_1_4_2 W_1_4_2_bar CIM_cell
X153 I143 O_1_4_3_3 WL_1_3 BL BLB W_1_4_3 W_1_4_3_bar CIM_cell
X154 I143 O_1_4_3_4 WL_1_3 BL BLB W_1_4_4 W_1_4_4_bar CIM_cell
X161 I144 O_1_4_4_1 WL_1_4 BL BLB W_1_4_1 W_1_4_1_bar CIM_cell
X162 I144 O_1_4_4_2 WL_1_4 BL BLB W_1_4_2 W_1_4_2_bar CIM_cell
X163 I144 O_1_4_4_3 WL_1_4 BL BLB W_1_4_3 W_1_4_3_bar CIM_cell
X164 I144 O_1_4_4_4 WL_1_4 BL BLB W_1_4_4 W_1_4_4_bar CIM_cell
X171 I151 O_1_5_1_1 WL_1_1 BL BLB W_1_5_1 W_1_5_1_bar CIM_cell
X172 I151 O_1_5_1_2 WL_1_1 BL BLB W_1_5_2 W_1_5_2_bar CIM_cell
X173 I151 O_1_5_1_3 WL_1_1 BL BLB W_1_5_3 W_1_5_3_bar CIM_cell
X174 I151 O_1_5_1_4 WL_1_1 BL BLB W_1_5_4 W_1_5_4_bar CIM_cell
X181 I152 O_1_5_2_1 WL_1_2 BL BLB W_1_5_1 W_1_5_1_bar CIM_cell
X182 I152 O_1_5_2_2 WL_1_2 BL BLB W_1_5_2 W_1_5_2_bar CIM_cell
X183 I152 O_1_5_2_3 WL_1_2 BL BLB W_1_5_3 W_1_5_3_bar CIM_cell
X184 I152 O_1_5_2_4 WL_1_2 BL BLB W_1_5_4 W_1_5_4_bar CIM_cell
X191 I153 O_1_5_3_1 WL_1_3 BL BLB W_1_5_1 W_1_5_1_bar CIM_cell
X192 I153 O_1_5_3_2 WL_1_3 BL BLB W_1_5_2 W_1_5_2_bar CIM_cell
X193 I153 O_1_5_3_3 WL_1_3 BL BLB W_1_5_3 W_1_5_3_bar CIM_cell
X194 I153 O_1_5_3_4 WL_1_3 BL BLB W_1_5_4 W_1_5_4_bar CIM_cell
X201 I154 O_1_5_4_1 WL_1_4 BL BLB W_1_5_1 W_1_5_1_bar CIM_cell
X202 I154 O_1_5_4_2 WL_1_4 BL BLB W_1_5_2 W_1_5_2_bar CIM_cell
X203 I154 O_1_5_4_3 WL_1_4 BL BLB W_1_5_3 W_1_5_3_bar CIM_cell
X204 I154 O_1_5_4_4 WL_1_4 BL BLB W_1_5_4 W_1_5_4_bar CIM_cell
X211 I161 O_1_6_1_1 WL_1_1 BL BLB W_1_6_1 W_1_6_1_bar CIM_cell
X212 I161 O_1_6_1_2 WL_1_1 BL BLB W_1_6_2 W_1_6_2_bar CIM_cell
X213 I161 O_1_6_1_3 WL_1_1 BL BLB W_1_6_3 W_1_6_3_bar CIM_cell
X214 I161 O_1_6_1_4 WL_1_1 BL BLB W_1_6_4 W_1_6_4_bar CIM_cell
X221 I162 O_1_6_2_1 WL_1_2 BL BLB W_1_6_1 W_1_6_1_bar CIM_cell
X222 I162 O_1_6_2_2 WL_1_2 BL BLB W_1_6_2 W_1_6_2_bar CIM_cell
X223 I162 O_1_6_2_3 WL_1_2 BL BLB W_1_6_3 W_1_6_3_bar CIM_cell
X224 I162 O_1_6_2_4 WL_1_2 BL BLB W_1_6_4 W_1_6_4_bar CIM_cell
X231 I163 O_1_6_3_1 WL_1_3 BL BLB W_1_6_1 W_1_6_1_bar CIM_cell
X232 I163 O_1_6_3_2 WL_1_3 BL BLB W_1_6_2 W_1_6_2_bar CIM_cell
X233 I163 O_1_6_3_3 WL_1_3 BL BLB W_1_6_3 W_1_6_3_bar CIM_cell
X234 I163 O_1_6_3_4 WL_1_3 BL BLB W_1_6_4 W_1_6_4_bar CIM_cell
X241 I164 O_1_6_4_1 WL_1_4 BL BLB W_1_6_1 W_1_6_1_bar CIM_cell
X242 I164 O_1_6_4_2 WL_1_4 BL BLB W_1_6_2 W_1_6_2_bar CIM_cell
X243 I164 O_1_6_4_3 WL_1_4 BL BLB W_1_6_3 W_1_6_3_bar CIM_cell
X244 I164 O_1_6_4_4 WL_1_4 BL BLB W_1_6_4 W_1_6_4_bar CIM_cell
X251 I171 O_1_7_1_1 WL_1_1 BL BLB W_1_7_1 W_1_7_1_bar CIM_cell
X252 I171 O_1_7_1_2 WL_1_1 BL BLB W_1_7_2 W_1_7_2_bar CIM_cell
X253 I171 O_1_7_1_3 WL_1_1 BL BLB W_1_7_3 W_1_7_3_bar CIM_cell
X254 I171 O_1_7_1_4 WL_1_1 BL BLB W_1_7_4 W_1_7_4_bar CIM_cell
X261 I172 O_1_7_2_1 WL_1_2 BL BLB W_1_7_1 W_1_7_1_bar CIM_cell
X262 I172 O_1_7_2_2 WL_1_2 BL BLB W_1_7_2 W_1_7_2_bar CIM_cell
X263 I172 O_1_7_2_3 WL_1_2 BL BLB W_1_7_3 W_1_7_3_bar CIM_cell
X264 I172 O_1_7_2_4 WL_1_2 BL BLB W_1_7_4 W_1_7_4_bar CIM_cell
X271 I173 O_1_7_3_1 WL_1_3 BL BLB W_1_7_1 W_1_7_1_bar CIM_cell
X272 I173 O_1_7_3_2 WL_1_3 BL BLB W_1_7_2 W_1_7_2_bar CIM_cell
X273 I173 O_1_7_3_3 WL_1_3 BL BLB W_1_7_3 W_1_7_3_bar CIM_cell
X274 I173 O_1_7_3_4 WL_1_3 BL BLB W_1_7_4 W_1_7_4_bar CIM_cell
X281 I174 O_1_7_4_1 WL_1_4 BL BLB W_1_7_1 W_1_7_1_bar CIM_cell
X282 I174 O_1_7_4_2 WL_1_4 BL BLB W_1_7_2 W_1_7_2_bar CIM_cell
X283 I174 O_1_7_4_3 WL_1_4 BL BLB W_1_7_3 W_1_7_3_bar CIM_cell
X284 I174 O_1_7_4_4 WL_1_4 BL BLB W_1_7_4 W_1_7_4_bar CIM_cell
X291 I181 O_1_8_1_1 WL_1_1 BL BLB W_1_8_1 W_1_8_1_bar CIM_cell
X292 I181 O_1_8_1_2 WL_1_1 BL BLB W_1_8_2 W_1_8_2_bar CIM_cell
X293 I181 O_1_8_1_3 WL_1_1 BL BLB W_1_8_3 W_1_8_3_bar CIM_cell
X294 I181 O_1_8_1_4 WL_1_1 BL BLB W_1_8_4 W_1_8_4_bar CIM_cell
X301 I182 O_1_8_2_1 WL_1_2 BL BLB W_1_8_1 W_1_8_1_bar CIM_cell
X302 I182 O_1_8_2_2 WL_1_2 BL BLB W_1_8_2 W_1_8_2_bar CIM_cell
X303 I182 O_1_8_2_3 WL_1_2 BL BLB W_1_8_3 W_1_8_3_bar CIM_cell
X304 I182 O_1_8_2_4 WL_1_2 BL BLB W_1_8_4 W_1_8_4_bar CIM_cell
X311 I183 O_1_8_3_1 WL_1_3 BL BLB W_1_8_1 W_1_8_1_bar CIM_cell
X312 I183 O_1_8_3_2 WL_1_3 BL BLB W_1_8_2 W_1_8_2_bar CIM_cell
X313 I183 O_1_8_3_3 WL_1_3 BL BLB W_1_8_3 W_1_8_3_bar CIM_cell
X314 I183 O_1_8_3_4 WL_1_3 BL BLB W_1_8_4 W_1_8_4_bar CIM_cell
X321 I184 O_1_8_4_1 WL_1_4 BL BLB W_1_8_1 W_1_8_1_bar CIM_cell
X322 I184 O_1_8_4_2 WL_1_4 BL BLB W_1_8_2 W_1_8_2_bar CIM_cell
X323 I184 O_1_8_4_3 WL_1_4 BL BLB W_1_8_3 W_1_8_3_bar CIM_cell
X324 I184 O_1_8_4_4 WL_1_4 BL BLB W_1_8_4 W_1_8_4_bar CIM_cell
X331 I191 O_1_9_1_1 WL_1_1 BL BLB W_1_9_1 W_1_9_1_bar CIM_cell
X332 I191 O_1_9_1_2 WL_1_1 BL BLB W_1_9_2 W_1_9_2_bar CIM_cell
X333 I191 O_1_9_1_3 WL_1_1 BL BLB W_1_9_3 W_1_9_3_bar CIM_cell
X334 I191 O_1_9_1_4 WL_1_1 BL BLB W_1_9_4 W_1_9_4_bar CIM_cell
X341 I192 O_1_9_2_1 WL_1_2 BL BLB W_1_9_1 W_1_9_1_bar CIM_cell
X342 I192 O_1_9_2_2 WL_1_2 BL BLB W_1_9_2 W_1_9_2_bar CIM_cell
X343 I192 O_1_9_2_3 WL_1_2 BL BLB W_1_9_3 W_1_9_3_bar CIM_cell
X344 I192 O_1_9_2_4 WL_1_2 BL BLB W_1_9_4 W_1_9_4_bar CIM_cell
X351 I193 O_1_9_3_1 WL_1_3 BL BLB W_1_9_1 W_1_9_1_bar CIM_cell
X352 I193 O_1_9_3_2 WL_1_3 BL BLB W_1_9_2 W_1_9_2_bar CIM_cell
X353 I193 O_1_9_3_3 WL_1_3 BL BLB W_1_9_3 W_1_9_3_bar CIM_cell
X354 I193 O_1_9_3_4 WL_1_3 BL BLB W_1_9_4 W_1_9_4_bar CIM_cell
X361 I194 O_1_9_4_1 WL_1_4 BL BLB W_1_9_1 W_1_9_1_bar CIM_cell
X362 I194 O_1_9_4_2 WL_1_4 BL BLB W_1_9_2 W_1_9_2_bar CIM_cell
X363 I194 O_1_9_4_3 WL_1_4 BL BLB W_1_9_3 W_1_9_3_bar CIM_cell
X364 I194 O_1_9_4_4 WL_1_4 BL BLB W_1_9_4 W_1_9_4_bar CIM_cell
X371 I1101 O_1_10_1_1 WL_1_1 BL BLB W_1_10_1 W_1_10_1_bar CIM_cell
X372 I1101 O_1_10_1_2 WL_1_1 BL BLB W_1_10_2 W_1_10_2_bar CIM_cell
X373 I1101 O_1_10_1_3 WL_1_1 BL BLB W_1_10_3 W_1_10_3_bar CIM_cell
X374 I1101 O_1_10_1_4 WL_1_1 BL BLB W_1_10_4 W_1_10_4_bar CIM_cell
X381 I1102 O_1_10_2_1 WL_1_2 BL BLB W_1_10_1 W_1_10_1_bar CIM_cell
X382 I1102 O_1_10_2_2 WL_1_2 BL BLB W_1_10_2 W_1_10_2_bar CIM_cell
X383 I1102 O_1_10_2_3 WL_1_2 BL BLB W_1_10_3 W_1_10_3_bar CIM_cell
X384 I1102 O_1_10_2_4 WL_1_2 BL BLB W_1_10_4 W_1_10_4_bar CIM_cell
X391 I1103 O_1_10_3_1 WL_1_3 BL BLB W_1_10_1 W_1_10_1_bar CIM_cell
X392 I1103 O_1_10_3_2 WL_1_3 BL BLB W_1_10_2 W_1_10_2_bar CIM_cell
X393 I1103 O_1_10_3_3 WL_1_3 BL BLB W_1_10_3 W_1_10_3_bar CIM_cell
X394 I1103 O_1_10_3_4 WL_1_3 BL BLB W_1_10_4 W_1_10_4_bar CIM_cell
X401 I1104 O_1_10_4_1 WL_1_4 BL BLB W_1_10_1 W_1_10_1_bar CIM_cell
X402 I1104 O_1_10_4_2 WL_1_4 BL BLB W_1_10_2 W_1_10_2_bar CIM_cell
X403 I1104 O_1_10_4_3 WL_1_4 BL BLB W_1_10_3 W_1_10_3_bar CIM_cell
X404 I1104 O_1_10_4_4 WL_1_4 BL BLB W_1_10_4 W_1_10_4_bar CIM_cell
X411 I1111 O_1_11_1_1 WL_1_1 BL BLB W_1_11_1 W_1_11_1_bar CIM_cell
X412 I1111 O_1_11_1_2 WL_1_1 BL BLB W_1_11_2 W_1_11_2_bar CIM_cell
X413 I1111 O_1_11_1_3 WL_1_1 BL BLB W_1_11_3 W_1_11_3_bar CIM_cell
X414 I1111 O_1_11_1_4 WL_1_1 BL BLB W_1_11_4 W_1_11_4_bar CIM_cell
X421 I1112 O_1_11_2_1 WL_1_2 BL BLB W_1_11_1 W_1_11_1_bar CIM_cell
X422 I1112 O_1_11_2_2 WL_1_2 BL BLB W_1_11_2 W_1_11_2_bar CIM_cell
X423 I1112 O_1_11_2_3 WL_1_2 BL BLB W_1_11_3 W_1_11_3_bar CIM_cell
X424 I1112 O_1_11_2_4 WL_1_2 BL BLB W_1_11_4 W_1_11_4_bar CIM_cell
X431 I1113 O_1_11_3_1 WL_1_3 BL BLB W_1_11_1 W_1_11_1_bar CIM_cell
X432 I1113 O_1_11_3_2 WL_1_3 BL BLB W_1_11_2 W_1_11_2_bar CIM_cell
X433 I1113 O_1_11_3_3 WL_1_3 BL BLB W_1_11_3 W_1_11_3_bar CIM_cell
X434 I1113 O_1_11_3_4 WL_1_3 BL BLB W_1_11_4 W_1_11_4_bar CIM_cell
X441 I1114 O_1_11_4_1 WL_1_4 BL BLB W_1_11_1 W_1_11_1_bar CIM_cell
X442 I1114 O_1_11_4_2 WL_1_4 BL BLB W_1_11_2 W_1_11_2_bar CIM_cell
X443 I1114 O_1_11_4_3 WL_1_4 BL BLB W_1_11_3 W_1_11_3_bar CIM_cell
X444 I1114 O_1_11_4_4 WL_1_4 BL BLB W_1_11_4 W_1_11_4_bar CIM_cell
X451 I1121 O_1_12_1_1 WL_1_1 BL BLB W_1_12_1 W_1_12_1_bar CIM_cell
X452 I1121 O_1_12_1_2 WL_1_1 BL BLB W_1_12_2 W_1_12_2_bar CIM_cell
X453 I1121 O_1_12_1_3 WL_1_1 BL BLB W_1_12_3 W_1_12_3_bar CIM_cell
X454 I1121 O_1_12_1_4 WL_1_1 BL BLB W_1_12_4 W_1_12_4_bar CIM_cell
X461 I1122 O_1_12_2_1 WL_1_2 BL BLB W_1_12_1 W_1_12_1_bar CIM_cell
X462 I1122 O_1_12_2_2 WL_1_2 BL BLB W_1_12_2 W_1_12_2_bar CIM_cell
X463 I1122 O_1_12_2_3 WL_1_2 BL BLB W_1_12_3 W_1_12_3_bar CIM_cell
X464 I1122 O_1_12_2_4 WL_1_2 BL BLB W_1_12_4 W_1_12_4_bar CIM_cell
X471 I1123 O_1_12_3_1 WL_1_3 BL BLB W_1_12_1 W_1_12_1_bar CIM_cell
X472 I1123 O_1_12_3_2 WL_1_3 BL BLB W_1_12_2 W_1_12_2_bar CIM_cell
X473 I1123 O_1_12_3_3 WL_1_3 BL BLB W_1_12_3 W_1_12_3_bar CIM_cell
X474 I1123 O_1_12_3_4 WL_1_3 BL BLB W_1_12_4 W_1_12_4_bar CIM_cell
X481 I1124 O_1_12_4_1 WL_1_4 BL BLB W_1_12_1 W_1_12_1_bar CIM_cell
X482 I1124 O_1_12_4_2 WL_1_4 BL BLB W_1_12_2 W_1_12_2_bar CIM_cell
X483 I1124 O_1_12_4_3 WL_1_4 BL BLB W_1_12_3 W_1_12_3_bar CIM_cell
X484 I1124 O_1_12_4_4 WL_1_4 BL BLB W_1_12_4 W_1_12_4_bar CIM_cell
X491 I1131 O_1_13_1_1 WL_1_1 BL BLB W_1_13_1 W_1_13_1_bar CIM_cell
X492 I1131 O_1_13_1_2 WL_1_1 BL BLB W_1_13_2 W_1_13_2_bar CIM_cell
X493 I1131 O_1_13_1_3 WL_1_1 BL BLB W_1_13_3 W_1_13_3_bar CIM_cell
X494 I1131 O_1_13_1_4 WL_1_1 BL BLB W_1_13_4 W_1_13_4_bar CIM_cell
X501 I1132 O_1_13_2_1 WL_1_2 BL BLB W_1_13_1 W_1_13_1_bar CIM_cell
X502 I1132 O_1_13_2_2 WL_1_2 BL BLB W_1_13_2 W_1_13_2_bar CIM_cell
X503 I1132 O_1_13_2_3 WL_1_2 BL BLB W_1_13_3 W_1_13_3_bar CIM_cell
X504 I1132 O_1_13_2_4 WL_1_2 BL BLB W_1_13_4 W_1_13_4_bar CIM_cell
X511 I1133 O_1_13_3_1 WL_1_3 BL BLB W_1_13_1 W_1_13_1_bar CIM_cell
X512 I1133 O_1_13_3_2 WL_1_3 BL BLB W_1_13_2 W_1_13_2_bar CIM_cell
X513 I1133 O_1_13_3_3 WL_1_3 BL BLB W_1_13_3 W_1_13_3_bar CIM_cell
X514 I1133 O_1_13_3_4 WL_1_3 BL BLB W_1_13_4 W_1_13_4_bar CIM_cell
X521 I1134 O_1_13_4_1 WL_1_4 BL BLB W_1_13_1 W_1_13_1_bar CIM_cell
X522 I1134 O_1_13_4_2 WL_1_4 BL BLB W_1_13_2 W_1_13_2_bar CIM_cell
X523 I1134 O_1_13_4_3 WL_1_4 BL BLB W_1_13_3 W_1_13_3_bar CIM_cell
X524 I1134 O_1_13_4_4 WL_1_4 BL BLB W_1_13_4 W_1_13_4_bar CIM_cell
X531 I1141 O_1_14_1_1 WL_1_1 BL BLB W_1_14_1 W_1_14_1_bar CIM_cell
X532 I1141 O_1_14_1_2 WL_1_1 BL BLB W_1_14_2 W_1_14_2_bar CIM_cell
X533 I1141 O_1_14_1_3 WL_1_1 BL BLB W_1_14_3 W_1_14_3_bar CIM_cell
X534 I1141 O_1_14_1_4 WL_1_1 BL BLB W_1_14_4 W_1_14_4_bar CIM_cell
X541 I1142 O_1_14_2_1 WL_1_2 BL BLB W_1_14_1 W_1_14_1_bar CIM_cell
X542 I1142 O_1_14_2_2 WL_1_2 BL BLB W_1_14_2 W_1_14_2_bar CIM_cell
X543 I1142 O_1_14_2_3 WL_1_2 BL BLB W_1_14_3 W_1_14_3_bar CIM_cell
X544 I1142 O_1_14_2_4 WL_1_2 BL BLB W_1_14_4 W_1_14_4_bar CIM_cell
X551 I1143 O_1_14_3_1 WL_1_3 BL BLB W_1_14_1 W_1_14_1_bar CIM_cell
X552 I1143 O_1_14_3_2 WL_1_3 BL BLB W_1_14_2 W_1_14_2_bar CIM_cell
X553 I1143 O_1_14_3_3 WL_1_3 BL BLB W_1_14_3 W_1_14_3_bar CIM_cell
X554 I1143 O_1_14_3_4 WL_1_3 BL BLB W_1_14_4 W_1_14_4_bar CIM_cell
X561 I1144 O_1_14_4_1 WL_1_4 BL BLB W_1_14_1 W_1_14_1_bar CIM_cell
X562 I1144 O_1_14_4_2 WL_1_4 BL BLB W_1_14_2 W_1_14_2_bar CIM_cell
X563 I1144 O_1_14_4_3 WL_1_4 BL BLB W_1_14_3 W_1_14_3_bar CIM_cell
X564 I1144 O_1_14_4_4 WL_1_4 BL BLB W_1_14_4 W_1_14_4_bar CIM_cell
X571 I1151 O_1_15_1_1 WL_1_1 BL BLB W_1_15_1 W_1_15_1_bar CIM_cell
X572 I1151 O_1_15_1_2 WL_1_1 BL BLB W_1_15_2 W_1_15_2_bar CIM_cell
X573 I1151 O_1_15_1_3 WL_1_1 BL BLB W_1_15_3 W_1_15_3_bar CIM_cell
X574 I1151 O_1_15_1_4 WL_1_1 BL BLB W_1_15_4 W_1_15_4_bar CIM_cell
X581 I1152 O_1_15_2_1 WL_1_2 BL BLB W_1_15_1 W_1_15_1_bar CIM_cell
X582 I1152 O_1_15_2_2 WL_1_2 BL BLB W_1_15_2 W_1_15_2_bar CIM_cell
X583 I1152 O_1_15_2_3 WL_1_2 BL BLB W_1_15_3 W_1_15_3_bar CIM_cell
X584 I1152 O_1_15_2_4 WL_1_2 BL BLB W_1_15_4 W_1_15_4_bar CIM_cell
X591 I1153 O_1_15_3_1 WL_1_3 BL BLB W_1_15_1 W_1_15_1_bar CIM_cell
X592 I1153 O_1_15_3_2 WL_1_3 BL BLB W_1_15_2 W_1_15_2_bar CIM_cell
X593 I1153 O_1_15_3_3 WL_1_3 BL BLB W_1_15_3 W_1_15_3_bar CIM_cell
X594 I1153 O_1_15_3_4 WL_1_3 BL BLB W_1_15_4 W_1_15_4_bar CIM_cell
X601 I1154 O_1_15_4_1 WL_1_4 BL BLB W_1_15_1 W_1_15_1_bar CIM_cell
X602 I1154 O_1_15_4_2 WL_1_4 BL BLB W_1_15_2 W_1_15_2_bar CIM_cell
X603 I1154 O_1_15_4_3 WL_1_4 BL BLB W_1_15_3 W_1_15_3_bar CIM_cell
X604 I1154 O_1_15_4_4 WL_1_4 BL BLB W_1_15_4 W_1_15_4_bar CIM_cell
X611 I1161 O_1_16_1_1 WL_1_1 BL BLB W_1_16_1 W_1_16_1_bar CIM_cell
X612 I1161 O_1_16_1_2 WL_1_1 BL BLB W_1_16_2 W_1_16_2_bar CIM_cell
X613 I1161 O_1_16_1_3 WL_1_1 BL BLB W_1_16_3 W_1_16_3_bar CIM_cell
X614 I1161 O_1_16_1_4 WL_1_1 BL BLB W_1_16_4 W_1_16_4_bar CIM_cell
X621 I1162 O_1_16_2_1 WL_1_2 BL BLB W_1_16_1 W_1_16_1_bar CIM_cell
X622 I1162 O_1_16_2_2 WL_1_2 BL BLB W_1_16_2 W_1_16_2_bar CIM_cell
X623 I1162 O_1_16_2_3 WL_1_2 BL BLB W_1_16_3 W_1_16_3_bar CIM_cell
X624 I1162 O_1_16_2_4 WL_1_2 BL BLB W_1_16_4 W_1_16_4_bar CIM_cell
X631 I1163 O_1_16_3_1 WL_1_3 BL BLB W_1_16_1 W_1_16_1_bar CIM_cell
X632 I1163 O_1_16_3_2 WL_1_3 BL BLB W_1_16_2 W_1_16_2_bar CIM_cell
X633 I1163 O_1_16_3_3 WL_1_3 BL BLB W_1_16_3 W_1_16_3_bar CIM_cell
X634 I1163 O_1_16_3_4 WL_1_3 BL BLB W_1_16_4 W_1_16_4_bar CIM_cell
X641 I1164 O_1_16_4_1 WL_1_4 BL BLB W_1_16_1 W_1_16_1_bar CIM_cell
X642 I1164 O_1_16_4_2 WL_1_4 BL BLB W_1_16_2 W_1_16_2_bar CIM_cell
X643 I1164 O_1_16_4_3 WL_1_4 BL BLB W_1_16_3 W_1_16_3_bar CIM_cell
X644 I1164 O_1_16_4_4 WL_1_4 BL BLB W_1_16_4 W_1_16_4_bar CIM_cell
X651 I1171 O_1_17_1_1 WL_1_1 BL BLB W_1_17_1 W_1_17_1_bar CIM_cell
X652 I1171 O_1_17_1_2 WL_1_1 BL BLB W_1_17_2 W_1_17_2_bar CIM_cell
X653 I1171 O_1_17_1_3 WL_1_1 BL BLB W_1_17_3 W_1_17_3_bar CIM_cell
X654 I1171 O_1_17_1_4 WL_1_1 BL BLB W_1_17_4 W_1_17_4_bar CIM_cell
X661 I1172 O_1_17_2_1 WL_1_2 BL BLB W_1_17_1 W_1_17_1_bar CIM_cell
X662 I1172 O_1_17_2_2 WL_1_2 BL BLB W_1_17_2 W_1_17_2_bar CIM_cell
X663 I1172 O_1_17_2_3 WL_1_2 BL BLB W_1_17_3 W_1_17_3_bar CIM_cell
X664 I1172 O_1_17_2_4 WL_1_2 BL BLB W_1_17_4 W_1_17_4_bar CIM_cell
X671 I1173 O_1_17_3_1 WL_1_3 BL BLB W_1_17_1 W_1_17_1_bar CIM_cell
X672 I1173 O_1_17_3_2 WL_1_3 BL BLB W_1_17_2 W_1_17_2_bar CIM_cell
X673 I1173 O_1_17_3_3 WL_1_3 BL BLB W_1_17_3 W_1_17_3_bar CIM_cell
X674 I1173 O_1_17_3_4 WL_1_3 BL BLB W_1_17_4 W_1_17_4_bar CIM_cell
X681 I1174 O_1_17_4_1 WL_1_4 BL BLB W_1_17_1 W_1_17_1_bar CIM_cell
X682 I1174 O_1_17_4_2 WL_1_4 BL BLB W_1_17_2 W_1_17_2_bar CIM_cell
X683 I1174 O_1_17_4_3 WL_1_4 BL BLB W_1_17_3 W_1_17_3_bar CIM_cell
X684 I1174 O_1_17_4_4 WL_1_4 BL BLB W_1_17_4 W_1_17_4_bar CIM_cell
X691 I1181 O_1_18_1_1 WL_1_1 BL BLB W_1_18_1 W_1_18_1_bar CIM_cell
X692 I1181 O_1_18_1_2 WL_1_1 BL BLB W_1_18_2 W_1_18_2_bar CIM_cell
X693 I1181 O_1_18_1_3 WL_1_1 BL BLB W_1_18_3 W_1_18_3_bar CIM_cell
X694 I1181 O_1_18_1_4 WL_1_1 BL BLB W_1_18_4 W_1_18_4_bar CIM_cell
X701 I1182 O_1_18_2_1 WL_1_2 BL BLB W_1_18_1 W_1_18_1_bar CIM_cell
X702 I1182 O_1_18_2_2 WL_1_2 BL BLB W_1_18_2 W_1_18_2_bar CIM_cell
X703 I1182 O_1_18_2_3 WL_1_2 BL BLB W_1_18_3 W_1_18_3_bar CIM_cell
X704 I1182 O_1_18_2_4 WL_1_2 BL BLB W_1_18_4 W_1_18_4_bar CIM_cell
X711 I1183 O_1_18_3_1 WL_1_3 BL BLB W_1_18_1 W_1_18_1_bar CIM_cell
X712 I1183 O_1_18_3_2 WL_1_3 BL BLB W_1_18_2 W_1_18_2_bar CIM_cell
X713 I1183 O_1_18_3_3 WL_1_3 BL BLB W_1_18_3 W_1_18_3_bar CIM_cell
X714 I1183 O_1_18_3_4 WL_1_3 BL BLB W_1_18_4 W_1_18_4_bar CIM_cell
X721 I1184 O_1_18_4_1 WL_1_4 BL BLB W_1_18_1 W_1_18_1_bar CIM_cell
X722 I1184 O_1_18_4_2 WL_1_4 BL BLB W_1_18_2 W_1_18_2_bar CIM_cell
X723 I1184 O_1_18_4_3 WL_1_4 BL BLB W_1_18_3 W_1_18_3_bar CIM_cell
X724 I1184 O_1_18_4_4 WL_1_4 BL BLB W_1_18_4 W_1_18_4_bar CIM_cell
X731 I1191 O_1_19_1_1 WL_1_1 BL BLB W_1_19_1 W_1_19_1_bar CIM_cell
X732 I1191 O_1_19_1_2 WL_1_1 BL BLB W_1_19_2 W_1_19_2_bar CIM_cell
X733 I1191 O_1_19_1_3 WL_1_1 BL BLB W_1_19_3 W_1_19_3_bar CIM_cell
X734 I1191 O_1_19_1_4 WL_1_1 BL BLB W_1_19_4 W_1_19_4_bar CIM_cell
X741 I1192 O_1_19_2_1 WL_1_2 BL BLB W_1_19_1 W_1_19_1_bar CIM_cell
X742 I1192 O_1_19_2_2 WL_1_2 BL BLB W_1_19_2 W_1_19_2_bar CIM_cell
X743 I1192 O_1_19_2_3 WL_1_2 BL BLB W_1_19_3 W_1_19_3_bar CIM_cell
X744 I1192 O_1_19_2_4 WL_1_2 BL BLB W_1_19_4 W_1_19_4_bar CIM_cell
X751 I1193 O_1_19_3_1 WL_1_3 BL BLB W_1_19_1 W_1_19_1_bar CIM_cell
X752 I1193 O_1_19_3_2 WL_1_3 BL BLB W_1_19_2 W_1_19_2_bar CIM_cell
X753 I1193 O_1_19_3_3 WL_1_3 BL BLB W_1_19_3 W_1_19_3_bar CIM_cell
X754 I1193 O_1_19_3_4 WL_1_3 BL BLB W_1_19_4 W_1_19_4_bar CIM_cell
X761 I1194 O_1_19_4_1 WL_1_4 BL BLB W_1_19_1 W_1_19_1_bar CIM_cell
X762 I1194 O_1_19_4_2 WL_1_4 BL BLB W_1_19_2 W_1_19_2_bar CIM_cell
X763 I1194 O_1_19_4_3 WL_1_4 BL BLB W_1_19_3 W_1_19_3_bar CIM_cell
X764 I1194 O_1_19_4_4 WL_1_4 BL BLB W_1_19_4 W_1_19_4_bar CIM_cell
X771 I1201 O_1_20_1_1 WL_1_1 BL BLB W_1_20_1 W_1_20_1_bar CIM_cell
X772 I1201 O_1_20_1_2 WL_1_1 BL BLB W_1_20_2 W_1_20_2_bar CIM_cell
X773 I1201 O_1_20_1_3 WL_1_1 BL BLB W_1_20_3 W_1_20_3_bar CIM_cell
X774 I1201 O_1_20_1_4 WL_1_1 BL BLB W_1_20_4 W_1_20_4_bar CIM_cell
X781 I1202 O_1_20_2_1 WL_1_2 BL BLB W_1_20_1 W_1_20_1_bar CIM_cell
X782 I1202 O_1_20_2_2 WL_1_2 BL BLB W_1_20_2 W_1_20_2_bar CIM_cell
X783 I1202 O_1_20_2_3 WL_1_2 BL BLB W_1_20_3 W_1_20_3_bar CIM_cell
X784 I1202 O_1_20_2_4 WL_1_2 BL BLB W_1_20_4 W_1_20_4_bar CIM_cell
X791 I1203 O_1_20_3_1 WL_1_3 BL BLB W_1_20_1 W_1_20_1_bar CIM_cell
X792 I1203 O_1_20_3_2 WL_1_3 BL BLB W_1_20_2 W_1_20_2_bar CIM_cell
X793 I1203 O_1_20_3_3 WL_1_3 BL BLB W_1_20_3 W_1_20_3_bar CIM_cell
X794 I1203 O_1_20_3_4 WL_1_3 BL BLB W_1_20_4 W_1_20_4_bar CIM_cell
X801 I1204 O_1_20_4_1 WL_1_4 BL BLB W_1_20_1 W_1_20_1_bar CIM_cell
X802 I1204 O_1_20_4_2 WL_1_4 BL BLB W_1_20_2 W_1_20_2_bar CIM_cell
X803 I1204 O_1_20_4_3 WL_1_4 BL BLB W_1_20_3 W_1_20_3_bar CIM_cell
X804 I1204 O_1_20_4_4 WL_1_4 BL BLB W_1_20_4 W_1_20_4_bar CIM_cell
X811 I1211 O_1_21_1_1 WL_1_1 BL BLB W_1_21_1 W_1_21_1_bar CIM_cell
X812 I1211 O_1_21_1_2 WL_1_1 BL BLB W_1_21_2 W_1_21_2_bar CIM_cell
X813 I1211 O_1_21_1_3 WL_1_1 BL BLB W_1_21_3 W_1_21_3_bar CIM_cell
X814 I1211 O_1_21_1_4 WL_1_1 BL BLB W_1_21_4 W_1_21_4_bar CIM_cell
X821 I1212 O_1_21_2_1 WL_1_2 BL BLB W_1_21_1 W_1_21_1_bar CIM_cell
X822 I1212 O_1_21_2_2 WL_1_2 BL BLB W_1_21_2 W_1_21_2_bar CIM_cell
X823 I1212 O_1_21_2_3 WL_1_2 BL BLB W_1_21_3 W_1_21_3_bar CIM_cell
X824 I1212 O_1_21_2_4 WL_1_2 BL BLB W_1_21_4 W_1_21_4_bar CIM_cell
X831 I1213 O_1_21_3_1 WL_1_3 BL BLB W_1_21_1 W_1_21_1_bar CIM_cell
X832 I1213 O_1_21_3_2 WL_1_3 BL BLB W_1_21_2 W_1_21_2_bar CIM_cell
X833 I1213 O_1_21_3_3 WL_1_3 BL BLB W_1_21_3 W_1_21_3_bar CIM_cell
X834 I1213 O_1_21_3_4 WL_1_3 BL BLB W_1_21_4 W_1_21_4_bar CIM_cell
X841 I1214 O_1_21_4_1 WL_1_4 BL BLB W_1_21_1 W_1_21_1_bar CIM_cell
X842 I1214 O_1_21_4_2 WL_1_4 BL BLB W_1_21_2 W_1_21_2_bar CIM_cell
X843 I1214 O_1_21_4_3 WL_1_4 BL BLB W_1_21_3 W_1_21_3_bar CIM_cell
X844 I1214 O_1_21_4_4 WL_1_4 BL BLB W_1_21_4 W_1_21_4_bar CIM_cell
X851 I1221 O_1_22_1_1 WL_1_1 BL BLB W_1_22_1 W_1_22_1_bar CIM_cell
X852 I1221 O_1_22_1_2 WL_1_1 BL BLB W_1_22_2 W_1_22_2_bar CIM_cell
X853 I1221 O_1_22_1_3 WL_1_1 BL BLB W_1_22_3 W_1_22_3_bar CIM_cell
X854 I1221 O_1_22_1_4 WL_1_1 BL BLB W_1_22_4 W_1_22_4_bar CIM_cell
X861 I1222 O_1_22_2_1 WL_1_2 BL BLB W_1_22_1 W_1_22_1_bar CIM_cell
X862 I1222 O_1_22_2_2 WL_1_2 BL BLB W_1_22_2 W_1_22_2_bar CIM_cell
X863 I1222 O_1_22_2_3 WL_1_2 BL BLB W_1_22_3 W_1_22_3_bar CIM_cell
X864 I1222 O_1_22_2_4 WL_1_2 BL BLB W_1_22_4 W_1_22_4_bar CIM_cell
X871 I1223 O_1_22_3_1 WL_1_3 BL BLB W_1_22_1 W_1_22_1_bar CIM_cell
X872 I1223 O_1_22_3_2 WL_1_3 BL BLB W_1_22_2 W_1_22_2_bar CIM_cell
X873 I1223 O_1_22_3_3 WL_1_3 BL BLB W_1_22_3 W_1_22_3_bar CIM_cell
X874 I1223 O_1_22_3_4 WL_1_3 BL BLB W_1_22_4 W_1_22_4_bar CIM_cell
X881 I1224 O_1_22_4_1 WL_1_4 BL BLB W_1_22_1 W_1_22_1_bar CIM_cell
X882 I1224 O_1_22_4_2 WL_1_4 BL BLB W_1_22_2 W_1_22_2_bar CIM_cell
X883 I1224 O_1_22_4_3 WL_1_4 BL BLB W_1_22_3 W_1_22_3_bar CIM_cell
X884 I1224 O_1_22_4_4 WL_1_4 BL BLB W_1_22_4 W_1_22_4_bar CIM_cell
X891 I1231 O_1_23_1_1 WL_1_1 BL BLB W_1_23_1 W_1_23_1_bar CIM_cell
X892 I1231 O_1_23_1_2 WL_1_1 BL BLB W_1_23_2 W_1_23_2_bar CIM_cell
X893 I1231 O_1_23_1_3 WL_1_1 BL BLB W_1_23_3 W_1_23_3_bar CIM_cell
X894 I1231 O_1_23_1_4 WL_1_1 BL BLB W_1_23_4 W_1_23_4_bar CIM_cell
X901 I1232 O_1_23_2_1 WL_1_2 BL BLB W_1_23_1 W_1_23_1_bar CIM_cell
X902 I1232 O_1_23_2_2 WL_1_2 BL BLB W_1_23_2 W_1_23_2_bar CIM_cell
X903 I1232 O_1_23_2_3 WL_1_2 BL BLB W_1_23_3 W_1_23_3_bar CIM_cell
X904 I1232 O_1_23_2_4 WL_1_2 BL BLB W_1_23_4 W_1_23_4_bar CIM_cell
X911 I1233 O_1_23_3_1 WL_1_3 BL BLB W_1_23_1 W_1_23_1_bar CIM_cell
X912 I1233 O_1_23_3_2 WL_1_3 BL BLB W_1_23_2 W_1_23_2_bar CIM_cell
X913 I1233 O_1_23_3_3 WL_1_3 BL BLB W_1_23_3 W_1_23_3_bar CIM_cell
X914 I1233 O_1_23_3_4 WL_1_3 BL BLB W_1_23_4 W_1_23_4_bar CIM_cell
X921 I1234 O_1_23_4_1 WL_1_4 BL BLB W_1_23_1 W_1_23_1_bar CIM_cell
X922 I1234 O_1_23_4_2 WL_1_4 BL BLB W_1_23_2 W_1_23_2_bar CIM_cell
X923 I1234 O_1_23_4_3 WL_1_4 BL BLB W_1_23_3 W_1_23_3_bar CIM_cell
X924 I1234 O_1_23_4_4 WL_1_4 BL BLB W_1_23_4 W_1_23_4_bar CIM_cell
X931 I1241 O_1_24_1_1 WL_1_1 BL BLB W_1_24_1 W_1_24_1_bar CIM_cell
X932 I1241 O_1_24_1_2 WL_1_1 BL BLB W_1_24_2 W_1_24_2_bar CIM_cell
X933 I1241 O_1_24_1_3 WL_1_1 BL BLB W_1_24_3 W_1_24_3_bar CIM_cell
X934 I1241 O_1_24_1_4 WL_1_1 BL BLB W_1_24_4 W_1_24_4_bar CIM_cell
X941 I1242 O_1_24_2_1 WL_1_2 BL BLB W_1_24_1 W_1_24_1_bar CIM_cell
X942 I1242 O_1_24_2_2 WL_1_2 BL BLB W_1_24_2 W_1_24_2_bar CIM_cell
X943 I1242 O_1_24_2_3 WL_1_2 BL BLB W_1_24_3 W_1_24_3_bar CIM_cell
X944 I1242 O_1_24_2_4 WL_1_2 BL BLB W_1_24_4 W_1_24_4_bar CIM_cell
X951 I1243 O_1_24_3_1 WL_1_3 BL BLB W_1_24_1 W_1_24_1_bar CIM_cell
X952 I1243 O_1_24_3_2 WL_1_3 BL BLB W_1_24_2 W_1_24_2_bar CIM_cell
X953 I1243 O_1_24_3_3 WL_1_3 BL BLB W_1_24_3 W_1_24_3_bar CIM_cell
X954 I1243 O_1_24_3_4 WL_1_3 BL BLB W_1_24_4 W_1_24_4_bar CIM_cell
X961 I1244 O_1_24_4_1 WL_1_4 BL BLB W_1_24_1 W_1_24_1_bar CIM_cell
X962 I1244 O_1_24_4_2 WL_1_4 BL BLB W_1_24_2 W_1_24_2_bar CIM_cell
X963 I1244 O_1_24_4_3 WL_1_4 BL BLB W_1_24_3 W_1_24_3_bar CIM_cell
X964 I1244 O_1_24_4_4 WL_1_4 BL BLB W_1_24_4 W_1_24_4_bar CIM_cell
X971 I1251 O_1_25_1_1 WL_1_1 BL BLB W_1_25_1 W_1_25_1_bar CIM_cell
X972 I1251 O_1_25_1_2 WL_1_1 BL BLB W_1_25_2 W_1_25_2_bar CIM_cell
X973 I1251 O_1_25_1_3 WL_1_1 BL BLB W_1_25_3 W_1_25_3_bar CIM_cell
X974 I1251 O_1_25_1_4 WL_1_1 BL BLB W_1_25_4 W_1_25_4_bar CIM_cell
X981 I1252 O_1_25_2_1 WL_1_2 BL BLB W_1_25_1 W_1_25_1_bar CIM_cell
X982 I1252 O_1_25_2_2 WL_1_2 BL BLB W_1_25_2 W_1_25_2_bar CIM_cell
X983 I1252 O_1_25_2_3 WL_1_2 BL BLB W_1_25_3 W_1_25_3_bar CIM_cell
X984 I1252 O_1_25_2_4 WL_1_2 BL BLB W_1_25_4 W_1_25_4_bar CIM_cell
X991 I1253 O_1_25_3_1 WL_1_3 BL BLB W_1_25_1 W_1_25_1_bar CIM_cell
X992 I1253 O_1_25_3_2 WL_1_3 BL BLB W_1_25_2 W_1_25_2_bar CIM_cell
X993 I1253 O_1_25_3_3 WL_1_3 BL BLB W_1_25_3 W_1_25_3_bar CIM_cell
X994 I1253 O_1_25_3_4 WL_1_3 BL BLB W_1_25_4 W_1_25_4_bar CIM_cell
X1001 I1254 O_1_25_4_1 WL_1_4 BL BLB W_1_25_1 W_1_25_1_bar CIM_cell
X1002 I1254 O_1_25_4_2 WL_1_4 BL BLB W_1_25_2 W_1_25_2_bar CIM_cell
X1003 I1254 O_1_25_4_3 WL_1_4 BL BLB W_1_25_3 W_1_25_3_bar CIM_cell
X1004 I1254 O_1_25_4_4 WL_1_4 BL BLB W_1_25_4 W_1_25_4_bar CIM_cell
X1011 I1261 O_1_26_1_1 WL_1_1 BL BLB W_1_26_1 W_1_26_1_bar CIM_cell
X1012 I1261 O_1_26_1_2 WL_1_1 BL BLB W_1_26_2 W_1_26_2_bar CIM_cell
X1013 I1261 O_1_26_1_3 WL_1_1 BL BLB W_1_26_3 W_1_26_3_bar CIM_cell
X1014 I1261 O_1_26_1_4 WL_1_1 BL BLB W_1_26_4 W_1_26_4_bar CIM_cell
X1021 I1262 O_1_26_2_1 WL_1_2 BL BLB W_1_26_1 W_1_26_1_bar CIM_cell
X1022 I1262 O_1_26_2_2 WL_1_2 BL BLB W_1_26_2 W_1_26_2_bar CIM_cell
X1023 I1262 O_1_26_2_3 WL_1_2 BL BLB W_1_26_3 W_1_26_3_bar CIM_cell
X1024 I1262 O_1_26_2_4 WL_1_2 BL BLB W_1_26_4 W_1_26_4_bar CIM_cell
X1031 I1263 O_1_26_3_1 WL_1_3 BL BLB W_1_26_1 W_1_26_1_bar CIM_cell
X1032 I1263 O_1_26_3_2 WL_1_3 BL BLB W_1_26_2 W_1_26_2_bar CIM_cell
X1033 I1263 O_1_26_3_3 WL_1_3 BL BLB W_1_26_3 W_1_26_3_bar CIM_cell
X1034 I1263 O_1_26_3_4 WL_1_3 BL BLB W_1_26_4 W_1_26_4_bar CIM_cell
X1041 I1264 O_1_26_4_1 WL_1_4 BL BLB W_1_26_1 W_1_26_1_bar CIM_cell
X1042 I1264 O_1_26_4_2 WL_1_4 BL BLB W_1_26_2 W_1_26_2_bar CIM_cell
X1043 I1264 O_1_26_4_3 WL_1_4 BL BLB W_1_26_3 W_1_26_3_bar CIM_cell
X1044 I1264 O_1_26_4_4 WL_1_4 BL BLB W_1_26_4 W_1_26_4_bar CIM_cell
X1051 I1271 O_1_27_1_1 WL_1_1 BL BLB W_1_27_1 W_1_27_1_bar CIM_cell
X1052 I1271 O_1_27_1_2 WL_1_1 BL BLB W_1_27_2 W_1_27_2_bar CIM_cell
X1053 I1271 O_1_27_1_3 WL_1_1 BL BLB W_1_27_3 W_1_27_3_bar CIM_cell
X1054 I1271 O_1_27_1_4 WL_1_1 BL BLB W_1_27_4 W_1_27_4_bar CIM_cell
X1061 I1272 O_1_27_2_1 WL_1_2 BL BLB W_1_27_1 W_1_27_1_bar CIM_cell
X1062 I1272 O_1_27_2_2 WL_1_2 BL BLB W_1_27_2 W_1_27_2_bar CIM_cell
X1063 I1272 O_1_27_2_3 WL_1_2 BL BLB W_1_27_3 W_1_27_3_bar CIM_cell
X1064 I1272 O_1_27_2_4 WL_1_2 BL BLB W_1_27_4 W_1_27_4_bar CIM_cell
X1071 I1273 O_1_27_3_1 WL_1_3 BL BLB W_1_27_1 W_1_27_1_bar CIM_cell
X1072 I1273 O_1_27_3_2 WL_1_3 BL BLB W_1_27_2 W_1_27_2_bar CIM_cell
X1073 I1273 O_1_27_3_3 WL_1_3 BL BLB W_1_27_3 W_1_27_3_bar CIM_cell
X1074 I1273 O_1_27_3_4 WL_1_3 BL BLB W_1_27_4 W_1_27_4_bar CIM_cell
X1081 I1274 O_1_27_4_1 WL_1_4 BL BLB W_1_27_1 W_1_27_1_bar CIM_cell
X1082 I1274 O_1_27_4_2 WL_1_4 BL BLB W_1_27_2 W_1_27_2_bar CIM_cell
X1083 I1274 O_1_27_4_3 WL_1_4 BL BLB W_1_27_3 W_1_27_3_bar CIM_cell
X1084 I1274 O_1_27_4_4 WL_1_4 BL BLB W_1_27_4 W_1_27_4_bar CIM_cell
X1091 I1281 O_1_28_1_1 WL_1_1 BL BLB W_1_28_1 W_1_28_1_bar CIM_cell
X1092 I1281 O_1_28_1_2 WL_1_1 BL BLB W_1_28_2 W_1_28_2_bar CIM_cell
X1093 I1281 O_1_28_1_3 WL_1_1 BL BLB W_1_28_3 W_1_28_3_bar CIM_cell
X1094 I1281 O_1_28_1_4 WL_1_1 BL BLB W_1_28_4 W_1_28_4_bar CIM_cell
X1101 I1282 O_1_28_2_1 WL_1_2 BL BLB W_1_28_1 W_1_28_1_bar CIM_cell
X1102 I1282 O_1_28_2_2 WL_1_2 BL BLB W_1_28_2 W_1_28_2_bar CIM_cell
X1103 I1282 O_1_28_2_3 WL_1_2 BL BLB W_1_28_3 W_1_28_3_bar CIM_cell
X1104 I1282 O_1_28_2_4 WL_1_2 BL BLB W_1_28_4 W_1_28_4_bar CIM_cell
X1111 I1283 O_1_28_3_1 WL_1_3 BL BLB W_1_28_1 W_1_28_1_bar CIM_cell
X1112 I1283 O_1_28_3_2 WL_1_3 BL BLB W_1_28_2 W_1_28_2_bar CIM_cell
X1113 I1283 O_1_28_3_3 WL_1_3 BL BLB W_1_28_3 W_1_28_3_bar CIM_cell
X1114 I1283 O_1_28_3_4 WL_1_3 BL BLB W_1_28_4 W_1_28_4_bar CIM_cell
X1121 I1284 O_1_28_4_1 WL_1_4 BL BLB W_1_28_1 W_1_28_1_bar CIM_cell
X1122 I1284 O_1_28_4_2 WL_1_4 BL BLB W_1_28_2 W_1_28_2_bar CIM_cell
X1123 I1284 O_1_28_4_3 WL_1_4 BL BLB W_1_28_3 W_1_28_3_bar CIM_cell
X1124 I1284 O_1_28_4_4 WL_1_4 BL BLB W_1_28_4 W_1_28_4_bar CIM_cell
X1131 I1291 O_1_29_1_1 WL_1_1 BL BLB W_1_29_1 W_1_29_1_bar CIM_cell
X1132 I1291 O_1_29_1_2 WL_1_1 BL BLB W_1_29_2 W_1_29_2_bar CIM_cell
X1133 I1291 O_1_29_1_3 WL_1_1 BL BLB W_1_29_3 W_1_29_3_bar CIM_cell
X1134 I1291 O_1_29_1_4 WL_1_1 BL BLB W_1_29_4 W_1_29_4_bar CIM_cell
X1141 I1292 O_1_29_2_1 WL_1_2 BL BLB W_1_29_1 W_1_29_1_bar CIM_cell
X1142 I1292 O_1_29_2_2 WL_1_2 BL BLB W_1_29_2 W_1_29_2_bar CIM_cell
X1143 I1292 O_1_29_2_3 WL_1_2 BL BLB W_1_29_3 W_1_29_3_bar CIM_cell
X1144 I1292 O_1_29_2_4 WL_1_2 BL BLB W_1_29_4 W_1_29_4_bar CIM_cell
X1151 I1293 O_1_29_3_1 WL_1_3 BL BLB W_1_29_1 W_1_29_1_bar CIM_cell
X1152 I1293 O_1_29_3_2 WL_1_3 BL BLB W_1_29_2 W_1_29_2_bar CIM_cell
X1153 I1293 O_1_29_3_3 WL_1_3 BL BLB W_1_29_3 W_1_29_3_bar CIM_cell
X1154 I1293 O_1_29_3_4 WL_1_3 BL BLB W_1_29_4 W_1_29_4_bar CIM_cell
X1161 I1294 O_1_29_4_1 WL_1_4 BL BLB W_1_29_1 W_1_29_1_bar CIM_cell
X1162 I1294 O_1_29_4_2 WL_1_4 BL BLB W_1_29_2 W_1_29_2_bar CIM_cell
X1163 I1294 O_1_29_4_3 WL_1_4 BL BLB W_1_29_3 W_1_29_3_bar CIM_cell
X1164 I1294 O_1_29_4_4 WL_1_4 BL BLB W_1_29_4 W_1_29_4_bar CIM_cell
X1171 I1301 O_1_30_1_1 WL_1_1 BL BLB W_1_30_1 W_1_30_1_bar CIM_cell
X1172 I1301 O_1_30_1_2 WL_1_1 BL BLB W_1_30_2 W_1_30_2_bar CIM_cell
X1173 I1301 O_1_30_1_3 WL_1_1 BL BLB W_1_30_3 W_1_30_3_bar CIM_cell
X1174 I1301 O_1_30_1_4 WL_1_1 BL BLB W_1_30_4 W_1_30_4_bar CIM_cell
X1181 I1302 O_1_30_2_1 WL_1_2 BL BLB W_1_30_1 W_1_30_1_bar CIM_cell
X1182 I1302 O_1_30_2_2 WL_1_2 BL BLB W_1_30_2 W_1_30_2_bar CIM_cell
X1183 I1302 O_1_30_2_3 WL_1_2 BL BLB W_1_30_3 W_1_30_3_bar CIM_cell
X1184 I1302 O_1_30_2_4 WL_1_2 BL BLB W_1_30_4 W_1_30_4_bar CIM_cell
X1191 I1303 O_1_30_3_1 WL_1_3 BL BLB W_1_30_1 W_1_30_1_bar CIM_cell
X1192 I1303 O_1_30_3_2 WL_1_3 BL BLB W_1_30_2 W_1_30_2_bar CIM_cell
X1193 I1303 O_1_30_3_3 WL_1_3 BL BLB W_1_30_3 W_1_30_3_bar CIM_cell
X1194 I1303 O_1_30_3_4 WL_1_3 BL BLB W_1_30_4 W_1_30_4_bar CIM_cell
X1201 I1304 O_1_30_4_1 WL_1_4 BL BLB W_1_30_1 W_1_30_1_bar CIM_cell
X1202 I1304 O_1_30_4_2 WL_1_4 BL BLB W_1_30_2 W_1_30_2_bar CIM_cell
X1203 I1304 O_1_30_4_3 WL_1_4 BL BLB W_1_30_3 W_1_30_3_bar CIM_cell
X1204 I1304 O_1_30_4_4 WL_1_4 BL BLB W_1_30_4 W_1_30_4_bar CIM_cell
X1211 I1311 O_1_31_1_1 WL_1_1 BL BLB W_1_31_1 W_1_31_1_bar CIM_cell
X1212 I1311 O_1_31_1_2 WL_1_1 BL BLB W_1_31_2 W_1_31_2_bar CIM_cell
X1213 I1311 O_1_31_1_3 WL_1_1 BL BLB W_1_31_3 W_1_31_3_bar CIM_cell
X1214 I1311 O_1_31_1_4 WL_1_1 BL BLB W_1_31_4 W_1_31_4_bar CIM_cell
X1221 I1312 O_1_31_2_1 WL_1_2 BL BLB W_1_31_1 W_1_31_1_bar CIM_cell
X1222 I1312 O_1_31_2_2 WL_1_2 BL BLB W_1_31_2 W_1_31_2_bar CIM_cell
X1223 I1312 O_1_31_2_3 WL_1_2 BL BLB W_1_31_3 W_1_31_3_bar CIM_cell
X1224 I1312 O_1_31_2_4 WL_1_2 BL BLB W_1_31_4 W_1_31_4_bar CIM_cell
X1231 I1313 O_1_31_3_1 WL_1_3 BL BLB W_1_31_1 W_1_31_1_bar CIM_cell
X1232 I1313 O_1_31_3_2 WL_1_3 BL BLB W_1_31_2 W_1_31_2_bar CIM_cell
X1233 I1313 O_1_31_3_3 WL_1_3 BL BLB W_1_31_3 W_1_31_3_bar CIM_cell
X1234 I1313 O_1_31_3_4 WL_1_3 BL BLB W_1_31_4 W_1_31_4_bar CIM_cell
X1241 I1314 O_1_31_4_1 WL_1_4 BL BLB W_1_31_1 W_1_31_1_bar CIM_cell
X1242 I1314 O_1_31_4_2 WL_1_4 BL BLB W_1_31_2 W_1_31_2_bar CIM_cell
X1243 I1314 O_1_31_4_3 WL_1_4 BL BLB W_1_31_3 W_1_31_3_bar CIM_cell
X1244 I1314 O_1_31_4_4 WL_1_4 BL BLB W_1_31_4 W_1_31_4_bar CIM_cell
X1251 I1321 O_1_32_1_1 WL_1_1 BL BLB W_1_32_1 W_1_32_1_bar CIM_cell
X1252 I1321 O_1_32_1_2 WL_1_1 BL BLB W_1_32_2 W_1_32_2_bar CIM_cell
X1253 I1321 O_1_32_1_3 WL_1_1 BL BLB W_1_32_3 W_1_32_3_bar CIM_cell
X1254 I1321 O_1_32_1_4 WL_1_1 BL BLB W_1_32_4 W_1_32_4_bar CIM_cell
X1261 I1322 O_1_32_2_1 WL_1_2 BL BLB W_1_32_1 W_1_32_1_bar CIM_cell
X1262 I1322 O_1_32_2_2 WL_1_2 BL BLB W_1_32_2 W_1_32_2_bar CIM_cell
X1263 I1322 O_1_32_2_3 WL_1_2 BL BLB W_1_32_3 W_1_32_3_bar CIM_cell
X1264 I1322 O_1_32_2_4 WL_1_2 BL BLB W_1_32_4 W_1_32_4_bar CIM_cell
X1271 I1323 O_1_32_3_1 WL_1_3 BL BLB W_1_32_1 W_1_32_1_bar CIM_cell
X1272 I1323 O_1_32_3_2 WL_1_3 BL BLB W_1_32_2 W_1_32_2_bar CIM_cell
X1273 I1323 O_1_32_3_3 WL_1_3 BL BLB W_1_32_3 W_1_32_3_bar CIM_cell
X1274 I1323 O_1_32_3_4 WL_1_3 BL BLB W_1_32_4 W_1_32_4_bar CIM_cell
X1281 I1324 O_1_32_4_1 WL_1_4 BL BLB W_1_32_1 W_1_32_1_bar CIM_cell
X1282 I1324 O_1_32_4_2 WL_1_4 BL BLB W_1_32_2 W_1_32_2_bar CIM_cell
X1283 I1324 O_1_32_4_3 WL_1_4 BL BLB W_1_32_3 W_1_32_3_bar CIM_cell
X1284 I1324 O_1_32_4_4 WL_1_4 BL BLB W_1_32_4 W_1_32_4_bar CIM_cell
X1291 I211 O_2_1_1_1 WL_2_1 BL BLB W_2_1_1 W_2_1_1_bar CIM_cell
X1292 I211 O_2_1_1_2 WL_2_1 BL BLB W_2_1_2 W_2_1_2_bar CIM_cell
X1293 I211 O_2_1_1_3 WL_2_1 BL BLB W_2_1_3 W_2_1_3_bar CIM_cell
X1294 I211 O_2_1_1_4 WL_2_1 BL BLB W_2_1_4 W_2_1_4_bar CIM_cell
X1301 I212 O_2_1_2_1 WL_2_2 BL BLB W_2_1_1 W_2_1_1_bar CIM_cell
X1302 I212 O_2_1_2_2 WL_2_2 BL BLB W_2_1_2 W_2_1_2_bar CIM_cell
X1303 I212 O_2_1_2_3 WL_2_2 BL BLB W_2_1_3 W_2_1_3_bar CIM_cell
X1304 I212 O_2_1_2_4 WL_2_2 BL BLB W_2_1_4 W_2_1_4_bar CIM_cell
X1311 I213 O_2_1_3_1 WL_2_3 BL BLB W_2_1_1 W_2_1_1_bar CIM_cell
X1312 I213 O_2_1_3_2 WL_2_3 BL BLB W_2_1_2 W_2_1_2_bar CIM_cell
X1313 I213 O_2_1_3_3 WL_2_3 BL BLB W_2_1_3 W_2_1_3_bar CIM_cell
X1314 I213 O_2_1_3_4 WL_2_3 BL BLB W_2_1_4 W_2_1_4_bar CIM_cell
X1321 I214 O_2_1_4_1 WL_2_4 BL BLB W_2_1_1 W_2_1_1_bar CIM_cell
X1322 I214 O_2_1_4_2 WL_2_4 BL BLB W_2_1_2 W_2_1_2_bar CIM_cell
X1323 I214 O_2_1_4_3 WL_2_4 BL BLB W_2_1_3 W_2_1_3_bar CIM_cell
X1324 I214 O_2_1_4_4 WL_2_4 BL BLB W_2_1_4 W_2_1_4_bar CIM_cell
X1331 I221 O_2_2_1_1 WL_2_1 BL BLB W_2_2_1 W_2_2_1_bar CIM_cell
X1332 I221 O_2_2_1_2 WL_2_1 BL BLB W_2_2_2 W_2_2_2_bar CIM_cell
X1333 I221 O_2_2_1_3 WL_2_1 BL BLB W_2_2_3 W_2_2_3_bar CIM_cell
X1334 I221 O_2_2_1_4 WL_2_1 BL BLB W_2_2_4 W_2_2_4_bar CIM_cell
X1341 I222 O_2_2_2_1 WL_2_2 BL BLB W_2_2_1 W_2_2_1_bar CIM_cell
X1342 I222 O_2_2_2_2 WL_2_2 BL BLB W_2_2_2 W_2_2_2_bar CIM_cell
X1343 I222 O_2_2_2_3 WL_2_2 BL BLB W_2_2_3 W_2_2_3_bar CIM_cell
X1344 I222 O_2_2_2_4 WL_2_2 BL BLB W_2_2_4 W_2_2_4_bar CIM_cell
X1351 I223 O_2_2_3_1 WL_2_3 BL BLB W_2_2_1 W_2_2_1_bar CIM_cell
X1352 I223 O_2_2_3_2 WL_2_3 BL BLB W_2_2_2 W_2_2_2_bar CIM_cell
X1353 I223 O_2_2_3_3 WL_2_3 BL BLB W_2_2_3 W_2_2_3_bar CIM_cell
X1354 I223 O_2_2_3_4 WL_2_3 BL BLB W_2_2_4 W_2_2_4_bar CIM_cell
X1361 I224 O_2_2_4_1 WL_2_4 BL BLB W_2_2_1 W_2_2_1_bar CIM_cell
X1362 I224 O_2_2_4_2 WL_2_4 BL BLB W_2_2_2 W_2_2_2_bar CIM_cell
X1363 I224 O_2_2_4_3 WL_2_4 BL BLB W_2_2_3 W_2_2_3_bar CIM_cell
X1364 I224 O_2_2_4_4 WL_2_4 BL BLB W_2_2_4 W_2_2_4_bar CIM_cell
X1371 I231 O_2_3_1_1 WL_2_1 BL BLB W_2_3_1 W_2_3_1_bar CIM_cell
X1372 I231 O_2_3_1_2 WL_2_1 BL BLB W_2_3_2 W_2_3_2_bar CIM_cell
X1373 I231 O_2_3_1_3 WL_2_1 BL BLB W_2_3_3 W_2_3_3_bar CIM_cell
X1374 I231 O_2_3_1_4 WL_2_1 BL BLB W_2_3_4 W_2_3_4_bar CIM_cell
X1381 I232 O_2_3_2_1 WL_2_2 BL BLB W_2_3_1 W_2_3_1_bar CIM_cell
X1382 I232 O_2_3_2_2 WL_2_2 BL BLB W_2_3_2 W_2_3_2_bar CIM_cell
X1383 I232 O_2_3_2_3 WL_2_2 BL BLB W_2_3_3 W_2_3_3_bar CIM_cell
X1384 I232 O_2_3_2_4 WL_2_2 BL BLB W_2_3_4 W_2_3_4_bar CIM_cell
X1391 I233 O_2_3_3_1 WL_2_3 BL BLB W_2_3_1 W_2_3_1_bar CIM_cell
X1392 I233 O_2_3_3_2 WL_2_3 BL BLB W_2_3_2 W_2_3_2_bar CIM_cell
X1393 I233 O_2_3_3_3 WL_2_3 BL BLB W_2_3_3 W_2_3_3_bar CIM_cell
X1394 I233 O_2_3_3_4 WL_2_3 BL BLB W_2_3_4 W_2_3_4_bar CIM_cell
X1401 I234 O_2_3_4_1 WL_2_4 BL BLB W_2_3_1 W_2_3_1_bar CIM_cell
X1402 I234 O_2_3_4_2 WL_2_4 BL BLB W_2_3_2 W_2_3_2_bar CIM_cell
X1403 I234 O_2_3_4_3 WL_2_4 BL BLB W_2_3_3 W_2_3_3_bar CIM_cell
X1404 I234 O_2_3_4_4 WL_2_4 BL BLB W_2_3_4 W_2_3_4_bar CIM_cell
X1411 I241 O_2_4_1_1 WL_2_1 BL BLB W_2_4_1 W_2_4_1_bar CIM_cell
X1412 I241 O_2_4_1_2 WL_2_1 BL BLB W_2_4_2 W_2_4_2_bar CIM_cell
X1413 I241 O_2_4_1_3 WL_2_1 BL BLB W_2_4_3 W_2_4_3_bar CIM_cell
X1414 I241 O_2_4_1_4 WL_2_1 BL BLB W_2_4_4 W_2_4_4_bar CIM_cell
X1421 I242 O_2_4_2_1 WL_2_2 BL BLB W_2_4_1 W_2_4_1_bar CIM_cell
X1422 I242 O_2_4_2_2 WL_2_2 BL BLB W_2_4_2 W_2_4_2_bar CIM_cell
X1423 I242 O_2_4_2_3 WL_2_2 BL BLB W_2_4_3 W_2_4_3_bar CIM_cell
X1424 I242 O_2_4_2_4 WL_2_2 BL BLB W_2_4_4 W_2_4_4_bar CIM_cell
X1431 I243 O_2_4_3_1 WL_2_3 BL BLB W_2_4_1 W_2_4_1_bar CIM_cell
X1432 I243 O_2_4_3_2 WL_2_3 BL BLB W_2_4_2 W_2_4_2_bar CIM_cell
X1433 I243 O_2_4_3_3 WL_2_3 BL BLB W_2_4_3 W_2_4_3_bar CIM_cell
X1434 I243 O_2_4_3_4 WL_2_3 BL BLB W_2_4_4 W_2_4_4_bar CIM_cell
X1441 I244 O_2_4_4_1 WL_2_4 BL BLB W_2_4_1 W_2_4_1_bar CIM_cell
X1442 I244 O_2_4_4_2 WL_2_4 BL BLB W_2_4_2 W_2_4_2_bar CIM_cell
X1443 I244 O_2_4_4_3 WL_2_4 BL BLB W_2_4_3 W_2_4_3_bar CIM_cell
X1444 I244 O_2_4_4_4 WL_2_4 BL BLB W_2_4_4 W_2_4_4_bar CIM_cell
X1451 I251 O_2_5_1_1 WL_2_1 BL BLB W_2_5_1 W_2_5_1_bar CIM_cell
X1452 I251 O_2_5_1_2 WL_2_1 BL BLB W_2_5_2 W_2_5_2_bar CIM_cell
X1453 I251 O_2_5_1_3 WL_2_1 BL BLB W_2_5_3 W_2_5_3_bar CIM_cell
X1454 I251 O_2_5_1_4 WL_2_1 BL BLB W_2_5_4 W_2_5_4_bar CIM_cell
X1461 I252 O_2_5_2_1 WL_2_2 BL BLB W_2_5_1 W_2_5_1_bar CIM_cell
X1462 I252 O_2_5_2_2 WL_2_2 BL BLB W_2_5_2 W_2_5_2_bar CIM_cell
X1463 I252 O_2_5_2_3 WL_2_2 BL BLB W_2_5_3 W_2_5_3_bar CIM_cell
X1464 I252 O_2_5_2_4 WL_2_2 BL BLB W_2_5_4 W_2_5_4_bar CIM_cell
X1471 I253 O_2_5_3_1 WL_2_3 BL BLB W_2_5_1 W_2_5_1_bar CIM_cell
X1472 I253 O_2_5_3_2 WL_2_3 BL BLB W_2_5_2 W_2_5_2_bar CIM_cell
X1473 I253 O_2_5_3_3 WL_2_3 BL BLB W_2_5_3 W_2_5_3_bar CIM_cell
X1474 I253 O_2_5_3_4 WL_2_3 BL BLB W_2_5_4 W_2_5_4_bar CIM_cell
X1481 I254 O_2_5_4_1 WL_2_4 BL BLB W_2_5_1 W_2_5_1_bar CIM_cell
X1482 I254 O_2_5_4_2 WL_2_4 BL BLB W_2_5_2 W_2_5_2_bar CIM_cell
X1483 I254 O_2_5_4_3 WL_2_4 BL BLB W_2_5_3 W_2_5_3_bar CIM_cell
X1484 I254 O_2_5_4_4 WL_2_4 BL BLB W_2_5_4 W_2_5_4_bar CIM_cell
X1491 I261 O_2_6_1_1 WL_2_1 BL BLB W_2_6_1 W_2_6_1_bar CIM_cell
X1492 I261 O_2_6_1_2 WL_2_1 BL BLB W_2_6_2 W_2_6_2_bar CIM_cell
X1493 I261 O_2_6_1_3 WL_2_1 BL BLB W_2_6_3 W_2_6_3_bar CIM_cell
X1494 I261 O_2_6_1_4 WL_2_1 BL BLB W_2_6_4 W_2_6_4_bar CIM_cell
X1501 I262 O_2_6_2_1 WL_2_2 BL BLB W_2_6_1 W_2_6_1_bar CIM_cell
X1502 I262 O_2_6_2_2 WL_2_2 BL BLB W_2_6_2 W_2_6_2_bar CIM_cell
X1503 I262 O_2_6_2_3 WL_2_2 BL BLB W_2_6_3 W_2_6_3_bar CIM_cell
X1504 I262 O_2_6_2_4 WL_2_2 BL BLB W_2_6_4 W_2_6_4_bar CIM_cell
X1511 I263 O_2_6_3_1 WL_2_3 BL BLB W_2_6_1 W_2_6_1_bar CIM_cell
X1512 I263 O_2_6_3_2 WL_2_3 BL BLB W_2_6_2 W_2_6_2_bar CIM_cell
X1513 I263 O_2_6_3_3 WL_2_3 BL BLB W_2_6_3 W_2_6_3_bar CIM_cell
X1514 I263 O_2_6_3_4 WL_2_3 BL BLB W_2_6_4 W_2_6_4_bar CIM_cell
X1521 I264 O_2_6_4_1 WL_2_4 BL BLB W_2_6_1 W_2_6_1_bar CIM_cell
X1522 I264 O_2_6_4_2 WL_2_4 BL BLB W_2_6_2 W_2_6_2_bar CIM_cell
X1523 I264 O_2_6_4_3 WL_2_4 BL BLB W_2_6_3 W_2_6_3_bar CIM_cell
X1524 I264 O_2_6_4_4 WL_2_4 BL BLB W_2_6_4 W_2_6_4_bar CIM_cell
X1531 I271 O_2_7_1_1 WL_2_1 BL BLB W_2_7_1 W_2_7_1_bar CIM_cell
X1532 I271 O_2_7_1_2 WL_2_1 BL BLB W_2_7_2 W_2_7_2_bar CIM_cell
X1533 I271 O_2_7_1_3 WL_2_1 BL BLB W_2_7_3 W_2_7_3_bar CIM_cell
X1534 I271 O_2_7_1_4 WL_2_1 BL BLB W_2_7_4 W_2_7_4_bar CIM_cell
X1541 I272 O_2_7_2_1 WL_2_2 BL BLB W_2_7_1 W_2_7_1_bar CIM_cell
X1542 I272 O_2_7_2_2 WL_2_2 BL BLB W_2_7_2 W_2_7_2_bar CIM_cell
X1543 I272 O_2_7_2_3 WL_2_2 BL BLB W_2_7_3 W_2_7_3_bar CIM_cell
X1544 I272 O_2_7_2_4 WL_2_2 BL BLB W_2_7_4 W_2_7_4_bar CIM_cell
X1551 I273 O_2_7_3_1 WL_2_3 BL BLB W_2_7_1 W_2_7_1_bar CIM_cell
X1552 I273 O_2_7_3_2 WL_2_3 BL BLB W_2_7_2 W_2_7_2_bar CIM_cell
X1553 I273 O_2_7_3_3 WL_2_3 BL BLB W_2_7_3 W_2_7_3_bar CIM_cell
X1554 I273 O_2_7_3_4 WL_2_3 BL BLB W_2_7_4 W_2_7_4_bar CIM_cell
X1561 I274 O_2_7_4_1 WL_2_4 BL BLB W_2_7_1 W_2_7_1_bar CIM_cell
X1562 I274 O_2_7_4_2 WL_2_4 BL BLB W_2_7_2 W_2_7_2_bar CIM_cell
X1563 I274 O_2_7_4_3 WL_2_4 BL BLB W_2_7_3 W_2_7_3_bar CIM_cell
X1564 I274 O_2_7_4_4 WL_2_4 BL BLB W_2_7_4 W_2_7_4_bar CIM_cell
X1571 I281 O_2_8_1_1 WL_2_1 BL BLB W_2_8_1 W_2_8_1_bar CIM_cell
X1572 I281 O_2_8_1_2 WL_2_1 BL BLB W_2_8_2 W_2_8_2_bar CIM_cell
X1573 I281 O_2_8_1_3 WL_2_1 BL BLB W_2_8_3 W_2_8_3_bar CIM_cell
X1574 I281 O_2_8_1_4 WL_2_1 BL BLB W_2_8_4 W_2_8_4_bar CIM_cell
X1581 I282 O_2_8_2_1 WL_2_2 BL BLB W_2_8_1 W_2_8_1_bar CIM_cell
X1582 I282 O_2_8_2_2 WL_2_2 BL BLB W_2_8_2 W_2_8_2_bar CIM_cell
X1583 I282 O_2_8_2_3 WL_2_2 BL BLB W_2_8_3 W_2_8_3_bar CIM_cell
X1584 I282 O_2_8_2_4 WL_2_2 BL BLB W_2_8_4 W_2_8_4_bar CIM_cell
X1591 I283 O_2_8_3_1 WL_2_3 BL BLB W_2_8_1 W_2_8_1_bar CIM_cell
X1592 I283 O_2_8_3_2 WL_2_3 BL BLB W_2_8_2 W_2_8_2_bar CIM_cell
X1593 I283 O_2_8_3_3 WL_2_3 BL BLB W_2_8_3 W_2_8_3_bar CIM_cell
X1594 I283 O_2_8_3_4 WL_2_3 BL BLB W_2_8_4 W_2_8_4_bar CIM_cell
X1601 I284 O_2_8_4_1 WL_2_4 BL BLB W_2_8_1 W_2_8_1_bar CIM_cell
X1602 I284 O_2_8_4_2 WL_2_4 BL BLB W_2_8_2 W_2_8_2_bar CIM_cell
X1603 I284 O_2_8_4_3 WL_2_4 BL BLB W_2_8_3 W_2_8_3_bar CIM_cell
X1604 I284 O_2_8_4_4 WL_2_4 BL BLB W_2_8_4 W_2_8_4_bar CIM_cell
X1611 I291 O_2_9_1_1 WL_2_1 BL BLB W_2_9_1 W_2_9_1_bar CIM_cell
X1612 I291 O_2_9_1_2 WL_2_1 BL BLB W_2_9_2 W_2_9_2_bar CIM_cell
X1613 I291 O_2_9_1_3 WL_2_1 BL BLB W_2_9_3 W_2_9_3_bar CIM_cell
X1614 I291 O_2_9_1_4 WL_2_1 BL BLB W_2_9_4 W_2_9_4_bar CIM_cell
X1621 I292 O_2_9_2_1 WL_2_2 BL BLB W_2_9_1 W_2_9_1_bar CIM_cell
X1622 I292 O_2_9_2_2 WL_2_2 BL BLB W_2_9_2 W_2_9_2_bar CIM_cell
X1623 I292 O_2_9_2_3 WL_2_2 BL BLB W_2_9_3 W_2_9_3_bar CIM_cell
X1624 I292 O_2_9_2_4 WL_2_2 BL BLB W_2_9_4 W_2_9_4_bar CIM_cell
X1631 I293 O_2_9_3_1 WL_2_3 BL BLB W_2_9_1 W_2_9_1_bar CIM_cell
X1632 I293 O_2_9_3_2 WL_2_3 BL BLB W_2_9_2 W_2_9_2_bar CIM_cell
X1633 I293 O_2_9_3_3 WL_2_3 BL BLB W_2_9_3 W_2_9_3_bar CIM_cell
X1634 I293 O_2_9_3_4 WL_2_3 BL BLB W_2_9_4 W_2_9_4_bar CIM_cell
X1641 I294 O_2_9_4_1 WL_2_4 BL BLB W_2_9_1 W_2_9_1_bar CIM_cell
X1642 I294 O_2_9_4_2 WL_2_4 BL BLB W_2_9_2 W_2_9_2_bar CIM_cell
X1643 I294 O_2_9_4_3 WL_2_4 BL BLB W_2_9_3 W_2_9_3_bar CIM_cell
X1644 I294 O_2_9_4_4 WL_2_4 BL BLB W_2_9_4 W_2_9_4_bar CIM_cell
X1651 I2101 O_2_10_1_1 WL_2_1 BL BLB W_2_10_1 W_2_10_1_bar CIM_cell
X1652 I2101 O_2_10_1_2 WL_2_1 BL BLB W_2_10_2 W_2_10_2_bar CIM_cell
X1653 I2101 O_2_10_1_3 WL_2_1 BL BLB W_2_10_3 W_2_10_3_bar CIM_cell
X1654 I2101 O_2_10_1_4 WL_2_1 BL BLB W_2_10_4 W_2_10_4_bar CIM_cell
X1661 I2102 O_2_10_2_1 WL_2_2 BL BLB W_2_10_1 W_2_10_1_bar CIM_cell
X1662 I2102 O_2_10_2_2 WL_2_2 BL BLB W_2_10_2 W_2_10_2_bar CIM_cell
X1663 I2102 O_2_10_2_3 WL_2_2 BL BLB W_2_10_3 W_2_10_3_bar CIM_cell
X1664 I2102 O_2_10_2_4 WL_2_2 BL BLB W_2_10_4 W_2_10_4_bar CIM_cell
X1671 I2103 O_2_10_3_1 WL_2_3 BL BLB W_2_10_1 W_2_10_1_bar CIM_cell
X1672 I2103 O_2_10_3_2 WL_2_3 BL BLB W_2_10_2 W_2_10_2_bar CIM_cell
X1673 I2103 O_2_10_3_3 WL_2_3 BL BLB W_2_10_3 W_2_10_3_bar CIM_cell
X1674 I2103 O_2_10_3_4 WL_2_3 BL BLB W_2_10_4 W_2_10_4_bar CIM_cell
X1681 I2104 O_2_10_4_1 WL_2_4 BL BLB W_2_10_1 W_2_10_1_bar CIM_cell
X1682 I2104 O_2_10_4_2 WL_2_4 BL BLB W_2_10_2 W_2_10_2_bar CIM_cell
X1683 I2104 O_2_10_4_3 WL_2_4 BL BLB W_2_10_3 W_2_10_3_bar CIM_cell
X1684 I2104 O_2_10_4_4 WL_2_4 BL BLB W_2_10_4 W_2_10_4_bar CIM_cell
X1691 I2111 O_2_11_1_1 WL_2_1 BL BLB W_2_11_1 W_2_11_1_bar CIM_cell
X1692 I2111 O_2_11_1_2 WL_2_1 BL BLB W_2_11_2 W_2_11_2_bar CIM_cell
X1693 I2111 O_2_11_1_3 WL_2_1 BL BLB W_2_11_3 W_2_11_3_bar CIM_cell
X1694 I2111 O_2_11_1_4 WL_2_1 BL BLB W_2_11_4 W_2_11_4_bar CIM_cell
X1701 I2112 O_2_11_2_1 WL_2_2 BL BLB W_2_11_1 W_2_11_1_bar CIM_cell
X1702 I2112 O_2_11_2_2 WL_2_2 BL BLB W_2_11_2 W_2_11_2_bar CIM_cell
X1703 I2112 O_2_11_2_3 WL_2_2 BL BLB W_2_11_3 W_2_11_3_bar CIM_cell
X1704 I2112 O_2_11_2_4 WL_2_2 BL BLB W_2_11_4 W_2_11_4_bar CIM_cell
X1711 I2113 O_2_11_3_1 WL_2_3 BL BLB W_2_11_1 W_2_11_1_bar CIM_cell
X1712 I2113 O_2_11_3_2 WL_2_3 BL BLB W_2_11_2 W_2_11_2_bar CIM_cell
X1713 I2113 O_2_11_3_3 WL_2_3 BL BLB W_2_11_3 W_2_11_3_bar CIM_cell
X1714 I2113 O_2_11_3_4 WL_2_3 BL BLB W_2_11_4 W_2_11_4_bar CIM_cell
X1721 I2114 O_2_11_4_1 WL_2_4 BL BLB W_2_11_1 W_2_11_1_bar CIM_cell
X1722 I2114 O_2_11_4_2 WL_2_4 BL BLB W_2_11_2 W_2_11_2_bar CIM_cell
X1723 I2114 O_2_11_4_3 WL_2_4 BL BLB W_2_11_3 W_2_11_3_bar CIM_cell
X1724 I2114 O_2_11_4_4 WL_2_4 BL BLB W_2_11_4 W_2_11_4_bar CIM_cell
X1731 I2121 O_2_12_1_1 WL_2_1 BL BLB W_2_12_1 W_2_12_1_bar CIM_cell
X1732 I2121 O_2_12_1_2 WL_2_1 BL BLB W_2_12_2 W_2_12_2_bar CIM_cell
X1733 I2121 O_2_12_1_3 WL_2_1 BL BLB W_2_12_3 W_2_12_3_bar CIM_cell
X1734 I2121 O_2_12_1_4 WL_2_1 BL BLB W_2_12_4 W_2_12_4_bar CIM_cell
X1741 I2122 O_2_12_2_1 WL_2_2 BL BLB W_2_12_1 W_2_12_1_bar CIM_cell
X1742 I2122 O_2_12_2_2 WL_2_2 BL BLB W_2_12_2 W_2_12_2_bar CIM_cell
X1743 I2122 O_2_12_2_3 WL_2_2 BL BLB W_2_12_3 W_2_12_3_bar CIM_cell
X1744 I2122 O_2_12_2_4 WL_2_2 BL BLB W_2_12_4 W_2_12_4_bar CIM_cell
X1751 I2123 O_2_12_3_1 WL_2_3 BL BLB W_2_12_1 W_2_12_1_bar CIM_cell
X1752 I2123 O_2_12_3_2 WL_2_3 BL BLB W_2_12_2 W_2_12_2_bar CIM_cell
X1753 I2123 O_2_12_3_3 WL_2_3 BL BLB W_2_12_3 W_2_12_3_bar CIM_cell
X1754 I2123 O_2_12_3_4 WL_2_3 BL BLB W_2_12_4 W_2_12_4_bar CIM_cell
X1761 I2124 O_2_12_4_1 WL_2_4 BL BLB W_2_12_1 W_2_12_1_bar CIM_cell
X1762 I2124 O_2_12_4_2 WL_2_4 BL BLB W_2_12_2 W_2_12_2_bar CIM_cell
X1763 I2124 O_2_12_4_3 WL_2_4 BL BLB W_2_12_3 W_2_12_3_bar CIM_cell
X1764 I2124 O_2_12_4_4 WL_2_4 BL BLB W_2_12_4 W_2_12_4_bar CIM_cell
X1771 I2131 O_2_13_1_1 WL_2_1 BL BLB W_2_13_1 W_2_13_1_bar CIM_cell
X1772 I2131 O_2_13_1_2 WL_2_1 BL BLB W_2_13_2 W_2_13_2_bar CIM_cell
X1773 I2131 O_2_13_1_3 WL_2_1 BL BLB W_2_13_3 W_2_13_3_bar CIM_cell
X1774 I2131 O_2_13_1_4 WL_2_1 BL BLB W_2_13_4 W_2_13_4_bar CIM_cell
X1781 I2132 O_2_13_2_1 WL_2_2 BL BLB W_2_13_1 W_2_13_1_bar CIM_cell
X1782 I2132 O_2_13_2_2 WL_2_2 BL BLB W_2_13_2 W_2_13_2_bar CIM_cell
X1783 I2132 O_2_13_2_3 WL_2_2 BL BLB W_2_13_3 W_2_13_3_bar CIM_cell
X1784 I2132 O_2_13_2_4 WL_2_2 BL BLB W_2_13_4 W_2_13_4_bar CIM_cell
X1791 I2133 O_2_13_3_1 WL_2_3 BL BLB W_2_13_1 W_2_13_1_bar CIM_cell
X1792 I2133 O_2_13_3_2 WL_2_3 BL BLB W_2_13_2 W_2_13_2_bar CIM_cell
X1793 I2133 O_2_13_3_3 WL_2_3 BL BLB W_2_13_3 W_2_13_3_bar CIM_cell
X1794 I2133 O_2_13_3_4 WL_2_3 BL BLB W_2_13_4 W_2_13_4_bar CIM_cell
X1801 I2134 O_2_13_4_1 WL_2_4 BL BLB W_2_13_1 W_2_13_1_bar CIM_cell
X1802 I2134 O_2_13_4_2 WL_2_4 BL BLB W_2_13_2 W_2_13_2_bar CIM_cell
X1803 I2134 O_2_13_4_3 WL_2_4 BL BLB W_2_13_3 W_2_13_3_bar CIM_cell
X1804 I2134 O_2_13_4_4 WL_2_4 BL BLB W_2_13_4 W_2_13_4_bar CIM_cell
X1811 I2141 O_2_14_1_1 WL_2_1 BL BLB W_2_14_1 W_2_14_1_bar CIM_cell
X1812 I2141 O_2_14_1_2 WL_2_1 BL BLB W_2_14_2 W_2_14_2_bar CIM_cell
X1813 I2141 O_2_14_1_3 WL_2_1 BL BLB W_2_14_3 W_2_14_3_bar CIM_cell
X1814 I2141 O_2_14_1_4 WL_2_1 BL BLB W_2_14_4 W_2_14_4_bar CIM_cell
X1821 I2142 O_2_14_2_1 WL_2_2 BL BLB W_2_14_1 W_2_14_1_bar CIM_cell
X1822 I2142 O_2_14_2_2 WL_2_2 BL BLB W_2_14_2 W_2_14_2_bar CIM_cell
X1823 I2142 O_2_14_2_3 WL_2_2 BL BLB W_2_14_3 W_2_14_3_bar CIM_cell
X1824 I2142 O_2_14_2_4 WL_2_2 BL BLB W_2_14_4 W_2_14_4_bar CIM_cell
X1831 I2143 O_2_14_3_1 WL_2_3 BL BLB W_2_14_1 W_2_14_1_bar CIM_cell
X1832 I2143 O_2_14_3_2 WL_2_3 BL BLB W_2_14_2 W_2_14_2_bar CIM_cell
X1833 I2143 O_2_14_3_3 WL_2_3 BL BLB W_2_14_3 W_2_14_3_bar CIM_cell
X1834 I2143 O_2_14_3_4 WL_2_3 BL BLB W_2_14_4 W_2_14_4_bar CIM_cell
X1841 I2144 O_2_14_4_1 WL_2_4 BL BLB W_2_14_1 W_2_14_1_bar CIM_cell
X1842 I2144 O_2_14_4_2 WL_2_4 BL BLB W_2_14_2 W_2_14_2_bar CIM_cell
X1843 I2144 O_2_14_4_3 WL_2_4 BL BLB W_2_14_3 W_2_14_3_bar CIM_cell
X1844 I2144 O_2_14_4_4 WL_2_4 BL BLB W_2_14_4 W_2_14_4_bar CIM_cell
X1851 I2151 O_2_15_1_1 WL_2_1 BL BLB W_2_15_1 W_2_15_1_bar CIM_cell
X1852 I2151 O_2_15_1_2 WL_2_1 BL BLB W_2_15_2 W_2_15_2_bar CIM_cell
X1853 I2151 O_2_15_1_3 WL_2_1 BL BLB W_2_15_3 W_2_15_3_bar CIM_cell
X1854 I2151 O_2_15_1_4 WL_2_1 BL BLB W_2_15_4 W_2_15_4_bar CIM_cell
X1861 I2152 O_2_15_2_1 WL_2_2 BL BLB W_2_15_1 W_2_15_1_bar CIM_cell
X1862 I2152 O_2_15_2_2 WL_2_2 BL BLB W_2_15_2 W_2_15_2_bar CIM_cell
X1863 I2152 O_2_15_2_3 WL_2_2 BL BLB W_2_15_3 W_2_15_3_bar CIM_cell
X1864 I2152 O_2_15_2_4 WL_2_2 BL BLB W_2_15_4 W_2_15_4_bar CIM_cell
X1871 I2153 O_2_15_3_1 WL_2_3 BL BLB W_2_15_1 W_2_15_1_bar CIM_cell
X1872 I2153 O_2_15_3_2 WL_2_3 BL BLB W_2_15_2 W_2_15_2_bar CIM_cell
X1873 I2153 O_2_15_3_3 WL_2_3 BL BLB W_2_15_3 W_2_15_3_bar CIM_cell
X1874 I2153 O_2_15_3_4 WL_2_3 BL BLB W_2_15_4 W_2_15_4_bar CIM_cell
X1881 I2154 O_2_15_4_1 WL_2_4 BL BLB W_2_15_1 W_2_15_1_bar CIM_cell
X1882 I2154 O_2_15_4_2 WL_2_4 BL BLB W_2_15_2 W_2_15_2_bar CIM_cell
X1883 I2154 O_2_15_4_3 WL_2_4 BL BLB W_2_15_3 W_2_15_3_bar CIM_cell
X1884 I2154 O_2_15_4_4 WL_2_4 BL BLB W_2_15_4 W_2_15_4_bar CIM_cell
X1891 I2161 O_2_16_1_1 WL_2_1 BL BLB W_2_16_1 W_2_16_1_bar CIM_cell
X1892 I2161 O_2_16_1_2 WL_2_1 BL BLB W_2_16_2 W_2_16_2_bar CIM_cell
X1893 I2161 O_2_16_1_3 WL_2_1 BL BLB W_2_16_3 W_2_16_3_bar CIM_cell
X1894 I2161 O_2_16_1_4 WL_2_1 BL BLB W_2_16_4 W_2_16_4_bar CIM_cell
X1901 I2162 O_2_16_2_1 WL_2_2 BL BLB W_2_16_1 W_2_16_1_bar CIM_cell
X1902 I2162 O_2_16_2_2 WL_2_2 BL BLB W_2_16_2 W_2_16_2_bar CIM_cell
X1903 I2162 O_2_16_2_3 WL_2_2 BL BLB W_2_16_3 W_2_16_3_bar CIM_cell
X1904 I2162 O_2_16_2_4 WL_2_2 BL BLB W_2_16_4 W_2_16_4_bar CIM_cell
X1911 I2163 O_2_16_3_1 WL_2_3 BL BLB W_2_16_1 W_2_16_1_bar CIM_cell
X1912 I2163 O_2_16_3_2 WL_2_3 BL BLB W_2_16_2 W_2_16_2_bar CIM_cell
X1913 I2163 O_2_16_3_3 WL_2_3 BL BLB W_2_16_3 W_2_16_3_bar CIM_cell
X1914 I2163 O_2_16_3_4 WL_2_3 BL BLB W_2_16_4 W_2_16_4_bar CIM_cell
X1921 I2164 O_2_16_4_1 WL_2_4 BL BLB W_2_16_1 W_2_16_1_bar CIM_cell
X1922 I2164 O_2_16_4_2 WL_2_4 BL BLB W_2_16_2 W_2_16_2_bar CIM_cell
X1923 I2164 O_2_16_4_3 WL_2_4 BL BLB W_2_16_3 W_2_16_3_bar CIM_cell
X1924 I2164 O_2_16_4_4 WL_2_4 BL BLB W_2_16_4 W_2_16_4_bar CIM_cell
X1931 I2171 O_2_17_1_1 WL_2_1 BL BLB W_2_17_1 W_2_17_1_bar CIM_cell
X1932 I2171 O_2_17_1_2 WL_2_1 BL BLB W_2_17_2 W_2_17_2_bar CIM_cell
X1933 I2171 O_2_17_1_3 WL_2_1 BL BLB W_2_17_3 W_2_17_3_bar CIM_cell
X1934 I2171 O_2_17_1_4 WL_2_1 BL BLB W_2_17_4 W_2_17_4_bar CIM_cell
X1941 I2172 O_2_17_2_1 WL_2_2 BL BLB W_2_17_1 W_2_17_1_bar CIM_cell
X1942 I2172 O_2_17_2_2 WL_2_2 BL BLB W_2_17_2 W_2_17_2_bar CIM_cell
X1943 I2172 O_2_17_2_3 WL_2_2 BL BLB W_2_17_3 W_2_17_3_bar CIM_cell
X1944 I2172 O_2_17_2_4 WL_2_2 BL BLB W_2_17_4 W_2_17_4_bar CIM_cell
X1951 I2173 O_2_17_3_1 WL_2_3 BL BLB W_2_17_1 W_2_17_1_bar CIM_cell
X1952 I2173 O_2_17_3_2 WL_2_3 BL BLB W_2_17_2 W_2_17_2_bar CIM_cell
X1953 I2173 O_2_17_3_3 WL_2_3 BL BLB W_2_17_3 W_2_17_3_bar CIM_cell
X1954 I2173 O_2_17_3_4 WL_2_3 BL BLB W_2_17_4 W_2_17_4_bar CIM_cell
X1961 I2174 O_2_17_4_1 WL_2_4 BL BLB W_2_17_1 W_2_17_1_bar CIM_cell
X1962 I2174 O_2_17_4_2 WL_2_4 BL BLB W_2_17_2 W_2_17_2_bar CIM_cell
X1963 I2174 O_2_17_4_3 WL_2_4 BL BLB W_2_17_3 W_2_17_3_bar CIM_cell
X1964 I2174 O_2_17_4_4 WL_2_4 BL BLB W_2_17_4 W_2_17_4_bar CIM_cell
X1971 I2181 O_2_18_1_1 WL_2_1 BL BLB W_2_18_1 W_2_18_1_bar CIM_cell
X1972 I2181 O_2_18_1_2 WL_2_1 BL BLB W_2_18_2 W_2_18_2_bar CIM_cell
X1973 I2181 O_2_18_1_3 WL_2_1 BL BLB W_2_18_3 W_2_18_3_bar CIM_cell
X1974 I2181 O_2_18_1_4 WL_2_1 BL BLB W_2_18_4 W_2_18_4_bar CIM_cell
X1981 I2182 O_2_18_2_1 WL_2_2 BL BLB W_2_18_1 W_2_18_1_bar CIM_cell
X1982 I2182 O_2_18_2_2 WL_2_2 BL BLB W_2_18_2 W_2_18_2_bar CIM_cell
X1983 I2182 O_2_18_2_3 WL_2_2 BL BLB W_2_18_3 W_2_18_3_bar CIM_cell
X1984 I2182 O_2_18_2_4 WL_2_2 BL BLB W_2_18_4 W_2_18_4_bar CIM_cell
X1991 I2183 O_2_18_3_1 WL_2_3 BL BLB W_2_18_1 W_2_18_1_bar CIM_cell
X1992 I2183 O_2_18_3_2 WL_2_3 BL BLB W_2_18_2 W_2_18_2_bar CIM_cell
X1993 I2183 O_2_18_3_3 WL_2_3 BL BLB W_2_18_3 W_2_18_3_bar CIM_cell
X1994 I2183 O_2_18_3_4 WL_2_3 BL BLB W_2_18_4 W_2_18_4_bar CIM_cell
X2001 I2184 O_2_18_4_1 WL_2_4 BL BLB W_2_18_1 W_2_18_1_bar CIM_cell
X2002 I2184 O_2_18_4_2 WL_2_4 BL BLB W_2_18_2 W_2_18_2_bar CIM_cell
X2003 I2184 O_2_18_4_3 WL_2_4 BL BLB W_2_18_3 W_2_18_3_bar CIM_cell
X2004 I2184 O_2_18_4_4 WL_2_4 BL BLB W_2_18_4 W_2_18_4_bar CIM_cell
X2011 I2191 O_2_19_1_1 WL_2_1 BL BLB W_2_19_1 W_2_19_1_bar CIM_cell
X2012 I2191 O_2_19_1_2 WL_2_1 BL BLB W_2_19_2 W_2_19_2_bar CIM_cell
X2013 I2191 O_2_19_1_3 WL_2_1 BL BLB W_2_19_3 W_2_19_3_bar CIM_cell
X2014 I2191 O_2_19_1_4 WL_2_1 BL BLB W_2_19_4 W_2_19_4_bar CIM_cell
X2021 I2192 O_2_19_2_1 WL_2_2 BL BLB W_2_19_1 W_2_19_1_bar CIM_cell
X2022 I2192 O_2_19_2_2 WL_2_2 BL BLB W_2_19_2 W_2_19_2_bar CIM_cell
X2023 I2192 O_2_19_2_3 WL_2_2 BL BLB W_2_19_3 W_2_19_3_bar CIM_cell
X2024 I2192 O_2_19_2_4 WL_2_2 BL BLB W_2_19_4 W_2_19_4_bar CIM_cell
X2031 I2193 O_2_19_3_1 WL_2_3 BL BLB W_2_19_1 W_2_19_1_bar CIM_cell
X2032 I2193 O_2_19_3_2 WL_2_3 BL BLB W_2_19_2 W_2_19_2_bar CIM_cell
X2033 I2193 O_2_19_3_3 WL_2_3 BL BLB W_2_19_3 W_2_19_3_bar CIM_cell
X2034 I2193 O_2_19_3_4 WL_2_3 BL BLB W_2_19_4 W_2_19_4_bar CIM_cell
X2041 I2194 O_2_19_4_1 WL_2_4 BL BLB W_2_19_1 W_2_19_1_bar CIM_cell
X2042 I2194 O_2_19_4_2 WL_2_4 BL BLB W_2_19_2 W_2_19_2_bar CIM_cell
X2043 I2194 O_2_19_4_3 WL_2_4 BL BLB W_2_19_3 W_2_19_3_bar CIM_cell
X2044 I2194 O_2_19_4_4 WL_2_4 BL BLB W_2_19_4 W_2_19_4_bar CIM_cell
X2051 I2201 O_2_20_1_1 WL_2_1 BL BLB W_2_20_1 W_2_20_1_bar CIM_cell
X2052 I2201 O_2_20_1_2 WL_2_1 BL BLB W_2_20_2 W_2_20_2_bar CIM_cell
X2053 I2201 O_2_20_1_3 WL_2_1 BL BLB W_2_20_3 W_2_20_3_bar CIM_cell
X2054 I2201 O_2_20_1_4 WL_2_1 BL BLB W_2_20_4 W_2_20_4_bar CIM_cell
X2061 I2202 O_2_20_2_1 WL_2_2 BL BLB W_2_20_1 W_2_20_1_bar CIM_cell
X2062 I2202 O_2_20_2_2 WL_2_2 BL BLB W_2_20_2 W_2_20_2_bar CIM_cell
X2063 I2202 O_2_20_2_3 WL_2_2 BL BLB W_2_20_3 W_2_20_3_bar CIM_cell
X2064 I2202 O_2_20_2_4 WL_2_2 BL BLB W_2_20_4 W_2_20_4_bar CIM_cell
X2071 I2203 O_2_20_3_1 WL_2_3 BL BLB W_2_20_1 W_2_20_1_bar CIM_cell
X2072 I2203 O_2_20_3_2 WL_2_3 BL BLB W_2_20_2 W_2_20_2_bar CIM_cell
X2073 I2203 O_2_20_3_3 WL_2_3 BL BLB W_2_20_3 W_2_20_3_bar CIM_cell
X2074 I2203 O_2_20_3_4 WL_2_3 BL BLB W_2_20_4 W_2_20_4_bar CIM_cell
X2081 I2204 O_2_20_4_1 WL_2_4 BL BLB W_2_20_1 W_2_20_1_bar CIM_cell
X2082 I2204 O_2_20_4_2 WL_2_4 BL BLB W_2_20_2 W_2_20_2_bar CIM_cell
X2083 I2204 O_2_20_4_3 WL_2_4 BL BLB W_2_20_3 W_2_20_3_bar CIM_cell
X2084 I2204 O_2_20_4_4 WL_2_4 BL BLB W_2_20_4 W_2_20_4_bar CIM_cell
X2091 I2211 O_2_21_1_1 WL_2_1 BL BLB W_2_21_1 W_2_21_1_bar CIM_cell
X2092 I2211 O_2_21_1_2 WL_2_1 BL BLB W_2_21_2 W_2_21_2_bar CIM_cell
X2093 I2211 O_2_21_1_3 WL_2_1 BL BLB W_2_21_3 W_2_21_3_bar CIM_cell
X2094 I2211 O_2_21_1_4 WL_2_1 BL BLB W_2_21_4 W_2_21_4_bar CIM_cell
X2101 I2212 O_2_21_2_1 WL_2_2 BL BLB W_2_21_1 W_2_21_1_bar CIM_cell
X2102 I2212 O_2_21_2_2 WL_2_2 BL BLB W_2_21_2 W_2_21_2_bar CIM_cell
X2103 I2212 O_2_21_2_3 WL_2_2 BL BLB W_2_21_3 W_2_21_3_bar CIM_cell
X2104 I2212 O_2_21_2_4 WL_2_2 BL BLB W_2_21_4 W_2_21_4_bar CIM_cell
X2111 I2213 O_2_21_3_1 WL_2_3 BL BLB W_2_21_1 W_2_21_1_bar CIM_cell
X2112 I2213 O_2_21_3_2 WL_2_3 BL BLB W_2_21_2 W_2_21_2_bar CIM_cell
X2113 I2213 O_2_21_3_3 WL_2_3 BL BLB W_2_21_3 W_2_21_3_bar CIM_cell
X2114 I2213 O_2_21_3_4 WL_2_3 BL BLB W_2_21_4 W_2_21_4_bar CIM_cell
X2121 I2214 O_2_21_4_1 WL_2_4 BL BLB W_2_21_1 W_2_21_1_bar CIM_cell
X2122 I2214 O_2_21_4_2 WL_2_4 BL BLB W_2_21_2 W_2_21_2_bar CIM_cell
X2123 I2214 O_2_21_4_3 WL_2_4 BL BLB W_2_21_3 W_2_21_3_bar CIM_cell
X2124 I2214 O_2_21_4_4 WL_2_4 BL BLB W_2_21_4 W_2_21_4_bar CIM_cell
X2131 I2221 O_2_22_1_1 WL_2_1 BL BLB W_2_22_1 W_2_22_1_bar CIM_cell
X2132 I2221 O_2_22_1_2 WL_2_1 BL BLB W_2_22_2 W_2_22_2_bar CIM_cell
X2133 I2221 O_2_22_1_3 WL_2_1 BL BLB W_2_22_3 W_2_22_3_bar CIM_cell
X2134 I2221 O_2_22_1_4 WL_2_1 BL BLB W_2_22_4 W_2_22_4_bar CIM_cell
X2141 I2222 O_2_22_2_1 WL_2_2 BL BLB W_2_22_1 W_2_22_1_bar CIM_cell
X2142 I2222 O_2_22_2_2 WL_2_2 BL BLB W_2_22_2 W_2_22_2_bar CIM_cell
X2143 I2222 O_2_22_2_3 WL_2_2 BL BLB W_2_22_3 W_2_22_3_bar CIM_cell
X2144 I2222 O_2_22_2_4 WL_2_2 BL BLB W_2_22_4 W_2_22_4_bar CIM_cell
X2151 I2223 O_2_22_3_1 WL_2_3 BL BLB W_2_22_1 W_2_22_1_bar CIM_cell
X2152 I2223 O_2_22_3_2 WL_2_3 BL BLB W_2_22_2 W_2_22_2_bar CIM_cell
X2153 I2223 O_2_22_3_3 WL_2_3 BL BLB W_2_22_3 W_2_22_3_bar CIM_cell
X2154 I2223 O_2_22_3_4 WL_2_3 BL BLB W_2_22_4 W_2_22_4_bar CIM_cell
X2161 I2224 O_2_22_4_1 WL_2_4 BL BLB W_2_22_1 W_2_22_1_bar CIM_cell
X2162 I2224 O_2_22_4_2 WL_2_4 BL BLB W_2_22_2 W_2_22_2_bar CIM_cell
X2163 I2224 O_2_22_4_3 WL_2_4 BL BLB W_2_22_3 W_2_22_3_bar CIM_cell
X2164 I2224 O_2_22_4_4 WL_2_4 BL BLB W_2_22_4 W_2_22_4_bar CIM_cell
X2171 I2231 O_2_23_1_1 WL_2_1 BL BLB W_2_23_1 W_2_23_1_bar CIM_cell
X2172 I2231 O_2_23_1_2 WL_2_1 BL BLB W_2_23_2 W_2_23_2_bar CIM_cell
X2173 I2231 O_2_23_1_3 WL_2_1 BL BLB W_2_23_3 W_2_23_3_bar CIM_cell
X2174 I2231 O_2_23_1_4 WL_2_1 BL BLB W_2_23_4 W_2_23_4_bar CIM_cell
X2181 I2232 O_2_23_2_1 WL_2_2 BL BLB W_2_23_1 W_2_23_1_bar CIM_cell
X2182 I2232 O_2_23_2_2 WL_2_2 BL BLB W_2_23_2 W_2_23_2_bar CIM_cell
X2183 I2232 O_2_23_2_3 WL_2_2 BL BLB W_2_23_3 W_2_23_3_bar CIM_cell
X2184 I2232 O_2_23_2_4 WL_2_2 BL BLB W_2_23_4 W_2_23_4_bar CIM_cell
X2191 I2233 O_2_23_3_1 WL_2_3 BL BLB W_2_23_1 W_2_23_1_bar CIM_cell
X2192 I2233 O_2_23_3_2 WL_2_3 BL BLB W_2_23_2 W_2_23_2_bar CIM_cell
X2193 I2233 O_2_23_3_3 WL_2_3 BL BLB W_2_23_3 W_2_23_3_bar CIM_cell
X2194 I2233 O_2_23_3_4 WL_2_3 BL BLB W_2_23_4 W_2_23_4_bar CIM_cell
X2201 I2234 O_2_23_4_1 WL_2_4 BL BLB W_2_23_1 W_2_23_1_bar CIM_cell
X2202 I2234 O_2_23_4_2 WL_2_4 BL BLB W_2_23_2 W_2_23_2_bar CIM_cell
X2203 I2234 O_2_23_4_3 WL_2_4 BL BLB W_2_23_3 W_2_23_3_bar CIM_cell
X2204 I2234 O_2_23_4_4 WL_2_4 BL BLB W_2_23_4 W_2_23_4_bar CIM_cell
X2211 I2241 O_2_24_1_1 WL_2_1 BL BLB W_2_24_1 W_2_24_1_bar CIM_cell
X2212 I2241 O_2_24_1_2 WL_2_1 BL BLB W_2_24_2 W_2_24_2_bar CIM_cell
X2213 I2241 O_2_24_1_3 WL_2_1 BL BLB W_2_24_3 W_2_24_3_bar CIM_cell
X2214 I2241 O_2_24_1_4 WL_2_1 BL BLB W_2_24_4 W_2_24_4_bar CIM_cell
X2221 I2242 O_2_24_2_1 WL_2_2 BL BLB W_2_24_1 W_2_24_1_bar CIM_cell
X2222 I2242 O_2_24_2_2 WL_2_2 BL BLB W_2_24_2 W_2_24_2_bar CIM_cell
X2223 I2242 O_2_24_2_3 WL_2_2 BL BLB W_2_24_3 W_2_24_3_bar CIM_cell
X2224 I2242 O_2_24_2_4 WL_2_2 BL BLB W_2_24_4 W_2_24_4_bar CIM_cell
X2231 I2243 O_2_24_3_1 WL_2_3 BL BLB W_2_24_1 W_2_24_1_bar CIM_cell
X2232 I2243 O_2_24_3_2 WL_2_3 BL BLB W_2_24_2 W_2_24_2_bar CIM_cell
X2233 I2243 O_2_24_3_3 WL_2_3 BL BLB W_2_24_3 W_2_24_3_bar CIM_cell
X2234 I2243 O_2_24_3_4 WL_2_3 BL BLB W_2_24_4 W_2_24_4_bar CIM_cell
X2241 I2244 O_2_24_4_1 WL_2_4 BL BLB W_2_24_1 W_2_24_1_bar CIM_cell
X2242 I2244 O_2_24_4_2 WL_2_4 BL BLB W_2_24_2 W_2_24_2_bar CIM_cell
X2243 I2244 O_2_24_4_3 WL_2_4 BL BLB W_2_24_3 W_2_24_3_bar CIM_cell
X2244 I2244 O_2_24_4_4 WL_2_4 BL BLB W_2_24_4 W_2_24_4_bar CIM_cell
X2251 I2251 O_2_25_1_1 WL_2_1 BL BLB W_2_25_1 W_2_25_1_bar CIM_cell
X2252 I2251 O_2_25_1_2 WL_2_1 BL BLB W_2_25_2 W_2_25_2_bar CIM_cell
X2253 I2251 O_2_25_1_3 WL_2_1 BL BLB W_2_25_3 W_2_25_3_bar CIM_cell
X2254 I2251 O_2_25_1_4 WL_2_1 BL BLB W_2_25_4 W_2_25_4_bar CIM_cell
X2261 I2252 O_2_25_2_1 WL_2_2 BL BLB W_2_25_1 W_2_25_1_bar CIM_cell
X2262 I2252 O_2_25_2_2 WL_2_2 BL BLB W_2_25_2 W_2_25_2_bar CIM_cell
X2263 I2252 O_2_25_2_3 WL_2_2 BL BLB W_2_25_3 W_2_25_3_bar CIM_cell
X2264 I2252 O_2_25_2_4 WL_2_2 BL BLB W_2_25_4 W_2_25_4_bar CIM_cell
X2271 I2253 O_2_25_3_1 WL_2_3 BL BLB W_2_25_1 W_2_25_1_bar CIM_cell
X2272 I2253 O_2_25_3_2 WL_2_3 BL BLB W_2_25_2 W_2_25_2_bar CIM_cell
X2273 I2253 O_2_25_3_3 WL_2_3 BL BLB W_2_25_3 W_2_25_3_bar CIM_cell
X2274 I2253 O_2_25_3_4 WL_2_3 BL BLB W_2_25_4 W_2_25_4_bar CIM_cell
X2281 I2254 O_2_25_4_1 WL_2_4 BL BLB W_2_25_1 W_2_25_1_bar CIM_cell
X2282 I2254 O_2_25_4_2 WL_2_4 BL BLB W_2_25_2 W_2_25_2_bar CIM_cell
X2283 I2254 O_2_25_4_3 WL_2_4 BL BLB W_2_25_3 W_2_25_3_bar CIM_cell
X2284 I2254 O_2_25_4_4 WL_2_4 BL BLB W_2_25_4 W_2_25_4_bar CIM_cell
X2291 I2261 O_2_26_1_1 WL_2_1 BL BLB W_2_26_1 W_2_26_1_bar CIM_cell
X2292 I2261 O_2_26_1_2 WL_2_1 BL BLB W_2_26_2 W_2_26_2_bar CIM_cell
X2293 I2261 O_2_26_1_3 WL_2_1 BL BLB W_2_26_3 W_2_26_3_bar CIM_cell
X2294 I2261 O_2_26_1_4 WL_2_1 BL BLB W_2_26_4 W_2_26_4_bar CIM_cell
X2301 I2262 O_2_26_2_1 WL_2_2 BL BLB W_2_26_1 W_2_26_1_bar CIM_cell
X2302 I2262 O_2_26_2_2 WL_2_2 BL BLB W_2_26_2 W_2_26_2_bar CIM_cell
X2303 I2262 O_2_26_2_3 WL_2_2 BL BLB W_2_26_3 W_2_26_3_bar CIM_cell
X2304 I2262 O_2_26_2_4 WL_2_2 BL BLB W_2_26_4 W_2_26_4_bar CIM_cell
X2311 I2263 O_2_26_3_1 WL_2_3 BL BLB W_2_26_1 W_2_26_1_bar CIM_cell
X2312 I2263 O_2_26_3_2 WL_2_3 BL BLB W_2_26_2 W_2_26_2_bar CIM_cell
X2313 I2263 O_2_26_3_3 WL_2_3 BL BLB W_2_26_3 W_2_26_3_bar CIM_cell
X2314 I2263 O_2_26_3_4 WL_2_3 BL BLB W_2_26_4 W_2_26_4_bar CIM_cell
X2321 I2264 O_2_26_4_1 WL_2_4 BL BLB W_2_26_1 W_2_26_1_bar CIM_cell
X2322 I2264 O_2_26_4_2 WL_2_4 BL BLB W_2_26_2 W_2_26_2_bar CIM_cell
X2323 I2264 O_2_26_4_3 WL_2_4 BL BLB W_2_26_3 W_2_26_3_bar CIM_cell
X2324 I2264 O_2_26_4_4 WL_2_4 BL BLB W_2_26_4 W_2_26_4_bar CIM_cell
X2331 I2271 O_2_27_1_1 WL_2_1 BL BLB W_2_27_1 W_2_27_1_bar CIM_cell
X2332 I2271 O_2_27_1_2 WL_2_1 BL BLB W_2_27_2 W_2_27_2_bar CIM_cell
X2333 I2271 O_2_27_1_3 WL_2_1 BL BLB W_2_27_3 W_2_27_3_bar CIM_cell
X2334 I2271 O_2_27_1_4 WL_2_1 BL BLB W_2_27_4 W_2_27_4_bar CIM_cell
X2341 I2272 O_2_27_2_1 WL_2_2 BL BLB W_2_27_1 W_2_27_1_bar CIM_cell
X2342 I2272 O_2_27_2_2 WL_2_2 BL BLB W_2_27_2 W_2_27_2_bar CIM_cell
X2343 I2272 O_2_27_2_3 WL_2_2 BL BLB W_2_27_3 W_2_27_3_bar CIM_cell
X2344 I2272 O_2_27_2_4 WL_2_2 BL BLB W_2_27_4 W_2_27_4_bar CIM_cell
X2351 I2273 O_2_27_3_1 WL_2_3 BL BLB W_2_27_1 W_2_27_1_bar CIM_cell
X2352 I2273 O_2_27_3_2 WL_2_3 BL BLB W_2_27_2 W_2_27_2_bar CIM_cell
X2353 I2273 O_2_27_3_3 WL_2_3 BL BLB W_2_27_3 W_2_27_3_bar CIM_cell
X2354 I2273 O_2_27_3_4 WL_2_3 BL BLB W_2_27_4 W_2_27_4_bar CIM_cell
X2361 I2274 O_2_27_4_1 WL_2_4 BL BLB W_2_27_1 W_2_27_1_bar CIM_cell
X2362 I2274 O_2_27_4_2 WL_2_4 BL BLB W_2_27_2 W_2_27_2_bar CIM_cell
X2363 I2274 O_2_27_4_3 WL_2_4 BL BLB W_2_27_3 W_2_27_3_bar CIM_cell
X2364 I2274 O_2_27_4_4 WL_2_4 BL BLB W_2_27_4 W_2_27_4_bar CIM_cell
X2371 I2281 O_2_28_1_1 WL_2_1 BL BLB W_2_28_1 W_2_28_1_bar CIM_cell
X2372 I2281 O_2_28_1_2 WL_2_1 BL BLB W_2_28_2 W_2_28_2_bar CIM_cell
X2373 I2281 O_2_28_1_3 WL_2_1 BL BLB W_2_28_3 W_2_28_3_bar CIM_cell
X2374 I2281 O_2_28_1_4 WL_2_1 BL BLB W_2_28_4 W_2_28_4_bar CIM_cell
X2381 I2282 O_2_28_2_1 WL_2_2 BL BLB W_2_28_1 W_2_28_1_bar CIM_cell
X2382 I2282 O_2_28_2_2 WL_2_2 BL BLB W_2_28_2 W_2_28_2_bar CIM_cell
X2383 I2282 O_2_28_2_3 WL_2_2 BL BLB W_2_28_3 W_2_28_3_bar CIM_cell
X2384 I2282 O_2_28_2_4 WL_2_2 BL BLB W_2_28_4 W_2_28_4_bar CIM_cell
X2391 I2283 O_2_28_3_1 WL_2_3 BL BLB W_2_28_1 W_2_28_1_bar CIM_cell
X2392 I2283 O_2_28_3_2 WL_2_3 BL BLB W_2_28_2 W_2_28_2_bar CIM_cell
X2393 I2283 O_2_28_3_3 WL_2_3 BL BLB W_2_28_3 W_2_28_3_bar CIM_cell
X2394 I2283 O_2_28_3_4 WL_2_3 BL BLB W_2_28_4 W_2_28_4_bar CIM_cell
X2401 I2284 O_2_28_4_1 WL_2_4 BL BLB W_2_28_1 W_2_28_1_bar CIM_cell
X2402 I2284 O_2_28_4_2 WL_2_4 BL BLB W_2_28_2 W_2_28_2_bar CIM_cell
X2403 I2284 O_2_28_4_3 WL_2_4 BL BLB W_2_28_3 W_2_28_3_bar CIM_cell
X2404 I2284 O_2_28_4_4 WL_2_4 BL BLB W_2_28_4 W_2_28_4_bar CIM_cell
X2411 I2291 O_2_29_1_1 WL_2_1 BL BLB W_2_29_1 W_2_29_1_bar CIM_cell
X2412 I2291 O_2_29_1_2 WL_2_1 BL BLB W_2_29_2 W_2_29_2_bar CIM_cell
X2413 I2291 O_2_29_1_3 WL_2_1 BL BLB W_2_29_3 W_2_29_3_bar CIM_cell
X2414 I2291 O_2_29_1_4 WL_2_1 BL BLB W_2_29_4 W_2_29_4_bar CIM_cell
X2421 I2292 O_2_29_2_1 WL_2_2 BL BLB W_2_29_1 W_2_29_1_bar CIM_cell
X2422 I2292 O_2_29_2_2 WL_2_2 BL BLB W_2_29_2 W_2_29_2_bar CIM_cell
X2423 I2292 O_2_29_2_3 WL_2_2 BL BLB W_2_29_3 W_2_29_3_bar CIM_cell
X2424 I2292 O_2_29_2_4 WL_2_2 BL BLB W_2_29_4 W_2_29_4_bar CIM_cell
X2431 I2293 O_2_29_3_1 WL_2_3 BL BLB W_2_29_1 W_2_29_1_bar CIM_cell
X2432 I2293 O_2_29_3_2 WL_2_3 BL BLB W_2_29_2 W_2_29_2_bar CIM_cell
X2433 I2293 O_2_29_3_3 WL_2_3 BL BLB W_2_29_3 W_2_29_3_bar CIM_cell
X2434 I2293 O_2_29_3_4 WL_2_3 BL BLB W_2_29_4 W_2_29_4_bar CIM_cell
X2441 I2294 O_2_29_4_1 WL_2_4 BL BLB W_2_29_1 W_2_29_1_bar CIM_cell
X2442 I2294 O_2_29_4_2 WL_2_4 BL BLB W_2_29_2 W_2_29_2_bar CIM_cell
X2443 I2294 O_2_29_4_3 WL_2_4 BL BLB W_2_29_3 W_2_29_3_bar CIM_cell
X2444 I2294 O_2_29_4_4 WL_2_4 BL BLB W_2_29_4 W_2_29_4_bar CIM_cell
X2451 I2301 O_2_30_1_1 WL_2_1 BL BLB W_2_30_1 W_2_30_1_bar CIM_cell
X2452 I2301 O_2_30_1_2 WL_2_1 BL BLB W_2_30_2 W_2_30_2_bar CIM_cell
X2453 I2301 O_2_30_1_3 WL_2_1 BL BLB W_2_30_3 W_2_30_3_bar CIM_cell
X2454 I2301 O_2_30_1_4 WL_2_1 BL BLB W_2_30_4 W_2_30_4_bar CIM_cell
X2461 I2302 O_2_30_2_1 WL_2_2 BL BLB W_2_30_1 W_2_30_1_bar CIM_cell
X2462 I2302 O_2_30_2_2 WL_2_2 BL BLB W_2_30_2 W_2_30_2_bar CIM_cell
X2463 I2302 O_2_30_2_3 WL_2_2 BL BLB W_2_30_3 W_2_30_3_bar CIM_cell
X2464 I2302 O_2_30_2_4 WL_2_2 BL BLB W_2_30_4 W_2_30_4_bar CIM_cell
X2471 I2303 O_2_30_3_1 WL_2_3 BL BLB W_2_30_1 W_2_30_1_bar CIM_cell
X2472 I2303 O_2_30_3_2 WL_2_3 BL BLB W_2_30_2 W_2_30_2_bar CIM_cell
X2473 I2303 O_2_30_3_3 WL_2_3 BL BLB W_2_30_3 W_2_30_3_bar CIM_cell
X2474 I2303 O_2_30_3_4 WL_2_3 BL BLB W_2_30_4 W_2_30_4_bar CIM_cell
X2481 I2304 O_2_30_4_1 WL_2_4 BL BLB W_2_30_1 W_2_30_1_bar CIM_cell
X2482 I2304 O_2_30_4_2 WL_2_4 BL BLB W_2_30_2 W_2_30_2_bar CIM_cell
X2483 I2304 O_2_30_4_3 WL_2_4 BL BLB W_2_30_3 W_2_30_3_bar CIM_cell
X2484 I2304 O_2_30_4_4 WL_2_4 BL BLB W_2_30_4 W_2_30_4_bar CIM_cell
X2491 I2311 O_2_31_1_1 WL_2_1 BL BLB W_2_31_1 W_2_31_1_bar CIM_cell
X2492 I2311 O_2_31_1_2 WL_2_1 BL BLB W_2_31_2 W_2_31_2_bar CIM_cell
X2493 I2311 O_2_31_1_3 WL_2_1 BL BLB W_2_31_3 W_2_31_3_bar CIM_cell
X2494 I2311 O_2_31_1_4 WL_2_1 BL BLB W_2_31_4 W_2_31_4_bar CIM_cell
X2501 I2312 O_2_31_2_1 WL_2_2 BL BLB W_2_31_1 W_2_31_1_bar CIM_cell
X2502 I2312 O_2_31_2_2 WL_2_2 BL BLB W_2_31_2 W_2_31_2_bar CIM_cell
X2503 I2312 O_2_31_2_3 WL_2_2 BL BLB W_2_31_3 W_2_31_3_bar CIM_cell
X2504 I2312 O_2_31_2_4 WL_2_2 BL BLB W_2_31_4 W_2_31_4_bar CIM_cell
X2511 I2313 O_2_31_3_1 WL_2_3 BL BLB W_2_31_1 W_2_31_1_bar CIM_cell
X2512 I2313 O_2_31_3_2 WL_2_3 BL BLB W_2_31_2 W_2_31_2_bar CIM_cell
X2513 I2313 O_2_31_3_3 WL_2_3 BL BLB W_2_31_3 W_2_31_3_bar CIM_cell
X2514 I2313 O_2_31_3_4 WL_2_3 BL BLB W_2_31_4 W_2_31_4_bar CIM_cell
X2521 I2314 O_2_31_4_1 WL_2_4 BL BLB W_2_31_1 W_2_31_1_bar CIM_cell
X2522 I2314 O_2_31_4_2 WL_2_4 BL BLB W_2_31_2 W_2_31_2_bar CIM_cell
X2523 I2314 O_2_31_4_3 WL_2_4 BL BLB W_2_31_3 W_2_31_3_bar CIM_cell
X2524 I2314 O_2_31_4_4 WL_2_4 BL BLB W_2_31_4 W_2_31_4_bar CIM_cell
X2531 I2321 O_2_32_1_1 WL_2_1 BL BLB W_2_32_1 W_2_32_1_bar CIM_cell
X2532 I2321 O_2_32_1_2 WL_2_1 BL BLB W_2_32_2 W_2_32_2_bar CIM_cell
X2533 I2321 O_2_32_1_3 WL_2_1 BL BLB W_2_32_3 W_2_32_3_bar CIM_cell
X2534 I2321 O_2_32_1_4 WL_2_1 BL BLB W_2_32_4 W_2_32_4_bar CIM_cell
X2541 I2322 O_2_32_2_1 WL_2_2 BL BLB W_2_32_1 W_2_32_1_bar CIM_cell
X2542 I2322 O_2_32_2_2 WL_2_2 BL BLB W_2_32_2 W_2_32_2_bar CIM_cell
X2543 I2322 O_2_32_2_3 WL_2_2 BL BLB W_2_32_3 W_2_32_3_bar CIM_cell
X2544 I2322 O_2_32_2_4 WL_2_2 BL BLB W_2_32_4 W_2_32_4_bar CIM_cell
X2551 I2323 O_2_32_3_1 WL_2_3 BL BLB W_2_32_1 W_2_32_1_bar CIM_cell
X2552 I2323 O_2_32_3_2 WL_2_3 BL BLB W_2_32_2 W_2_32_2_bar CIM_cell
X2553 I2323 O_2_32_3_3 WL_2_3 BL BLB W_2_32_3 W_2_32_3_bar CIM_cell
X2554 I2323 O_2_32_3_4 WL_2_3 BL BLB W_2_32_4 W_2_32_4_bar CIM_cell
X2561 I2324 O_2_32_4_1 WL_2_4 BL BLB W_2_32_1 W_2_32_1_bar CIM_cell
X2562 I2324 O_2_32_4_2 WL_2_4 BL BLB W_2_32_2 W_2_32_2_bar CIM_cell
X2563 I2324 O_2_32_4_3 WL_2_4 BL BLB W_2_32_3 W_2_32_3_bar CIM_cell
X2564 I2324 O_2_32_4_4 WL_2_4 BL BLB W_2_32_4 W_2_32_4_bar CIM_cell
X2571 I311 O_3_1_1_1 WL_3_1 BL BLB W_3_1_1 W_3_1_1_bar CIM_cell
X2572 I311 O_3_1_1_2 WL_3_1 BL BLB W_3_1_2 W_3_1_2_bar CIM_cell
X2573 I311 O_3_1_1_3 WL_3_1 BL BLB W_3_1_3 W_3_1_3_bar CIM_cell
X2574 I311 O_3_1_1_4 WL_3_1 BL BLB W_3_1_4 W_3_1_4_bar CIM_cell
X2581 I312 O_3_1_2_1 WL_3_2 BL BLB W_3_1_1 W_3_1_1_bar CIM_cell
X2582 I312 O_3_1_2_2 WL_3_2 BL BLB W_3_1_2 W_3_1_2_bar CIM_cell
X2583 I312 O_3_1_2_3 WL_3_2 BL BLB W_3_1_3 W_3_1_3_bar CIM_cell
X2584 I312 O_3_1_2_4 WL_3_2 BL BLB W_3_1_4 W_3_1_4_bar CIM_cell
X2591 I313 O_3_1_3_1 WL_3_3 BL BLB W_3_1_1 W_3_1_1_bar CIM_cell
X2592 I313 O_3_1_3_2 WL_3_3 BL BLB W_3_1_2 W_3_1_2_bar CIM_cell
X2593 I313 O_3_1_3_3 WL_3_3 BL BLB W_3_1_3 W_3_1_3_bar CIM_cell
X2594 I313 O_3_1_3_4 WL_3_3 BL BLB W_3_1_4 W_3_1_4_bar CIM_cell
X2601 I314 O_3_1_4_1 WL_3_4 BL BLB W_3_1_1 W_3_1_1_bar CIM_cell
X2602 I314 O_3_1_4_2 WL_3_4 BL BLB W_3_1_2 W_3_1_2_bar CIM_cell
X2603 I314 O_3_1_4_3 WL_3_4 BL BLB W_3_1_3 W_3_1_3_bar CIM_cell
X2604 I314 O_3_1_4_4 WL_3_4 BL BLB W_3_1_4 W_3_1_4_bar CIM_cell
X2611 I321 O_3_2_1_1 WL_3_1 BL BLB W_3_2_1 W_3_2_1_bar CIM_cell
X2612 I321 O_3_2_1_2 WL_3_1 BL BLB W_3_2_2 W_3_2_2_bar CIM_cell
X2613 I321 O_3_2_1_3 WL_3_1 BL BLB W_3_2_3 W_3_2_3_bar CIM_cell
X2614 I321 O_3_2_1_4 WL_3_1 BL BLB W_3_2_4 W_3_2_4_bar CIM_cell
X2621 I322 O_3_2_2_1 WL_3_2 BL BLB W_3_2_1 W_3_2_1_bar CIM_cell
X2622 I322 O_3_2_2_2 WL_3_2 BL BLB W_3_2_2 W_3_2_2_bar CIM_cell
X2623 I322 O_3_2_2_3 WL_3_2 BL BLB W_3_2_3 W_3_2_3_bar CIM_cell
X2624 I322 O_3_2_2_4 WL_3_2 BL BLB W_3_2_4 W_3_2_4_bar CIM_cell
X2631 I323 O_3_2_3_1 WL_3_3 BL BLB W_3_2_1 W_3_2_1_bar CIM_cell
X2632 I323 O_3_2_3_2 WL_3_3 BL BLB W_3_2_2 W_3_2_2_bar CIM_cell
X2633 I323 O_3_2_3_3 WL_3_3 BL BLB W_3_2_3 W_3_2_3_bar CIM_cell
X2634 I323 O_3_2_3_4 WL_3_3 BL BLB W_3_2_4 W_3_2_4_bar CIM_cell
X2641 I324 O_3_2_4_1 WL_3_4 BL BLB W_3_2_1 W_3_2_1_bar CIM_cell
X2642 I324 O_3_2_4_2 WL_3_4 BL BLB W_3_2_2 W_3_2_2_bar CIM_cell
X2643 I324 O_3_2_4_3 WL_3_4 BL BLB W_3_2_3 W_3_2_3_bar CIM_cell
X2644 I324 O_3_2_4_4 WL_3_4 BL BLB W_3_2_4 W_3_2_4_bar CIM_cell
X2651 I331 O_3_3_1_1 WL_3_1 BL BLB W_3_3_1 W_3_3_1_bar CIM_cell
X2652 I331 O_3_3_1_2 WL_3_1 BL BLB W_3_3_2 W_3_3_2_bar CIM_cell
X2653 I331 O_3_3_1_3 WL_3_1 BL BLB W_3_3_3 W_3_3_3_bar CIM_cell
X2654 I331 O_3_3_1_4 WL_3_1 BL BLB W_3_3_4 W_3_3_4_bar CIM_cell
X2661 I332 O_3_3_2_1 WL_3_2 BL BLB W_3_3_1 W_3_3_1_bar CIM_cell
X2662 I332 O_3_3_2_2 WL_3_2 BL BLB W_3_3_2 W_3_3_2_bar CIM_cell
X2663 I332 O_3_3_2_3 WL_3_2 BL BLB W_3_3_3 W_3_3_3_bar CIM_cell
X2664 I332 O_3_3_2_4 WL_3_2 BL BLB W_3_3_4 W_3_3_4_bar CIM_cell
X2671 I333 O_3_3_3_1 WL_3_3 BL BLB W_3_3_1 W_3_3_1_bar CIM_cell
X2672 I333 O_3_3_3_2 WL_3_3 BL BLB W_3_3_2 W_3_3_2_bar CIM_cell
X2673 I333 O_3_3_3_3 WL_3_3 BL BLB W_3_3_3 W_3_3_3_bar CIM_cell
X2674 I333 O_3_3_3_4 WL_3_3 BL BLB W_3_3_4 W_3_3_4_bar CIM_cell
X2681 I334 O_3_3_4_1 WL_3_4 BL BLB W_3_3_1 W_3_3_1_bar CIM_cell
X2682 I334 O_3_3_4_2 WL_3_4 BL BLB W_3_3_2 W_3_3_2_bar CIM_cell
X2683 I334 O_3_3_4_3 WL_3_4 BL BLB W_3_3_3 W_3_3_3_bar CIM_cell
X2684 I334 O_3_3_4_4 WL_3_4 BL BLB W_3_3_4 W_3_3_4_bar CIM_cell
X2691 I341 O_3_4_1_1 WL_3_1 BL BLB W_3_4_1 W_3_4_1_bar CIM_cell
X2692 I341 O_3_4_1_2 WL_3_1 BL BLB W_3_4_2 W_3_4_2_bar CIM_cell
X2693 I341 O_3_4_1_3 WL_3_1 BL BLB W_3_4_3 W_3_4_3_bar CIM_cell
X2694 I341 O_3_4_1_4 WL_3_1 BL BLB W_3_4_4 W_3_4_4_bar CIM_cell
X2701 I342 O_3_4_2_1 WL_3_2 BL BLB W_3_4_1 W_3_4_1_bar CIM_cell
X2702 I342 O_3_4_2_2 WL_3_2 BL BLB W_3_4_2 W_3_4_2_bar CIM_cell
X2703 I342 O_3_4_2_3 WL_3_2 BL BLB W_3_4_3 W_3_4_3_bar CIM_cell
X2704 I342 O_3_4_2_4 WL_3_2 BL BLB W_3_4_4 W_3_4_4_bar CIM_cell
X2711 I343 O_3_4_3_1 WL_3_3 BL BLB W_3_4_1 W_3_4_1_bar CIM_cell
X2712 I343 O_3_4_3_2 WL_3_3 BL BLB W_3_4_2 W_3_4_2_bar CIM_cell
X2713 I343 O_3_4_3_3 WL_3_3 BL BLB W_3_4_3 W_3_4_3_bar CIM_cell
X2714 I343 O_3_4_3_4 WL_3_3 BL BLB W_3_4_4 W_3_4_4_bar CIM_cell
X2721 I344 O_3_4_4_1 WL_3_4 BL BLB W_3_4_1 W_3_4_1_bar CIM_cell
X2722 I344 O_3_4_4_2 WL_3_4 BL BLB W_3_4_2 W_3_4_2_bar CIM_cell
X2723 I344 O_3_4_4_3 WL_3_4 BL BLB W_3_4_3 W_3_4_3_bar CIM_cell
X2724 I344 O_3_4_4_4 WL_3_4 BL BLB W_3_4_4 W_3_4_4_bar CIM_cell
X2731 I351 O_3_5_1_1 WL_3_1 BL BLB W_3_5_1 W_3_5_1_bar CIM_cell
X2732 I351 O_3_5_1_2 WL_3_1 BL BLB W_3_5_2 W_3_5_2_bar CIM_cell
X2733 I351 O_3_5_1_3 WL_3_1 BL BLB W_3_5_3 W_3_5_3_bar CIM_cell
X2734 I351 O_3_5_1_4 WL_3_1 BL BLB W_3_5_4 W_3_5_4_bar CIM_cell
X2741 I352 O_3_5_2_1 WL_3_2 BL BLB W_3_5_1 W_3_5_1_bar CIM_cell
X2742 I352 O_3_5_2_2 WL_3_2 BL BLB W_3_5_2 W_3_5_2_bar CIM_cell
X2743 I352 O_3_5_2_3 WL_3_2 BL BLB W_3_5_3 W_3_5_3_bar CIM_cell
X2744 I352 O_3_5_2_4 WL_3_2 BL BLB W_3_5_4 W_3_5_4_bar CIM_cell
X2751 I353 O_3_5_3_1 WL_3_3 BL BLB W_3_5_1 W_3_5_1_bar CIM_cell
X2752 I353 O_3_5_3_2 WL_3_3 BL BLB W_3_5_2 W_3_5_2_bar CIM_cell
X2753 I353 O_3_5_3_3 WL_3_3 BL BLB W_3_5_3 W_3_5_3_bar CIM_cell
X2754 I353 O_3_5_3_4 WL_3_3 BL BLB W_3_5_4 W_3_5_4_bar CIM_cell
X2761 I354 O_3_5_4_1 WL_3_4 BL BLB W_3_5_1 W_3_5_1_bar CIM_cell
X2762 I354 O_3_5_4_2 WL_3_4 BL BLB W_3_5_2 W_3_5_2_bar CIM_cell
X2763 I354 O_3_5_4_3 WL_3_4 BL BLB W_3_5_3 W_3_5_3_bar CIM_cell
X2764 I354 O_3_5_4_4 WL_3_4 BL BLB W_3_5_4 W_3_5_4_bar CIM_cell
X2771 I361 O_3_6_1_1 WL_3_1 BL BLB W_3_6_1 W_3_6_1_bar CIM_cell
X2772 I361 O_3_6_1_2 WL_3_1 BL BLB W_3_6_2 W_3_6_2_bar CIM_cell
X2773 I361 O_3_6_1_3 WL_3_1 BL BLB W_3_6_3 W_3_6_3_bar CIM_cell
X2774 I361 O_3_6_1_4 WL_3_1 BL BLB W_3_6_4 W_3_6_4_bar CIM_cell
X2781 I362 O_3_6_2_1 WL_3_2 BL BLB W_3_6_1 W_3_6_1_bar CIM_cell
X2782 I362 O_3_6_2_2 WL_3_2 BL BLB W_3_6_2 W_3_6_2_bar CIM_cell
X2783 I362 O_3_6_2_3 WL_3_2 BL BLB W_3_6_3 W_3_6_3_bar CIM_cell
X2784 I362 O_3_6_2_4 WL_3_2 BL BLB W_3_6_4 W_3_6_4_bar CIM_cell
X2791 I363 O_3_6_3_1 WL_3_3 BL BLB W_3_6_1 W_3_6_1_bar CIM_cell
X2792 I363 O_3_6_3_2 WL_3_3 BL BLB W_3_6_2 W_3_6_2_bar CIM_cell
X2793 I363 O_3_6_3_3 WL_3_3 BL BLB W_3_6_3 W_3_6_3_bar CIM_cell
X2794 I363 O_3_6_3_4 WL_3_3 BL BLB W_3_6_4 W_3_6_4_bar CIM_cell
X2801 I364 O_3_6_4_1 WL_3_4 BL BLB W_3_6_1 W_3_6_1_bar CIM_cell
X2802 I364 O_3_6_4_2 WL_3_4 BL BLB W_3_6_2 W_3_6_2_bar CIM_cell
X2803 I364 O_3_6_4_3 WL_3_4 BL BLB W_3_6_3 W_3_6_3_bar CIM_cell
X2804 I364 O_3_6_4_4 WL_3_4 BL BLB W_3_6_4 W_3_6_4_bar CIM_cell
X2811 I371 O_3_7_1_1 WL_3_1 BL BLB W_3_7_1 W_3_7_1_bar CIM_cell
X2812 I371 O_3_7_1_2 WL_3_1 BL BLB W_3_7_2 W_3_7_2_bar CIM_cell
X2813 I371 O_3_7_1_3 WL_3_1 BL BLB W_3_7_3 W_3_7_3_bar CIM_cell
X2814 I371 O_3_7_1_4 WL_3_1 BL BLB W_3_7_4 W_3_7_4_bar CIM_cell
X2821 I372 O_3_7_2_1 WL_3_2 BL BLB W_3_7_1 W_3_7_1_bar CIM_cell
X2822 I372 O_3_7_2_2 WL_3_2 BL BLB W_3_7_2 W_3_7_2_bar CIM_cell
X2823 I372 O_3_7_2_3 WL_3_2 BL BLB W_3_7_3 W_3_7_3_bar CIM_cell
X2824 I372 O_3_7_2_4 WL_3_2 BL BLB W_3_7_4 W_3_7_4_bar CIM_cell
X2831 I373 O_3_7_3_1 WL_3_3 BL BLB W_3_7_1 W_3_7_1_bar CIM_cell
X2832 I373 O_3_7_3_2 WL_3_3 BL BLB W_3_7_2 W_3_7_2_bar CIM_cell
X2833 I373 O_3_7_3_3 WL_3_3 BL BLB W_3_7_3 W_3_7_3_bar CIM_cell
X2834 I373 O_3_7_3_4 WL_3_3 BL BLB W_3_7_4 W_3_7_4_bar CIM_cell
X2841 I374 O_3_7_4_1 WL_3_4 BL BLB W_3_7_1 W_3_7_1_bar CIM_cell
X2842 I374 O_3_7_4_2 WL_3_4 BL BLB W_3_7_2 W_3_7_2_bar CIM_cell
X2843 I374 O_3_7_4_3 WL_3_4 BL BLB W_3_7_3 W_3_7_3_bar CIM_cell
X2844 I374 O_3_7_4_4 WL_3_4 BL BLB W_3_7_4 W_3_7_4_bar CIM_cell
X2851 I381 O_3_8_1_1 WL_3_1 BL BLB W_3_8_1 W_3_8_1_bar CIM_cell
X2852 I381 O_3_8_1_2 WL_3_1 BL BLB W_3_8_2 W_3_8_2_bar CIM_cell
X2853 I381 O_3_8_1_3 WL_3_1 BL BLB W_3_8_3 W_3_8_3_bar CIM_cell
X2854 I381 O_3_8_1_4 WL_3_1 BL BLB W_3_8_4 W_3_8_4_bar CIM_cell
X2861 I382 O_3_8_2_1 WL_3_2 BL BLB W_3_8_1 W_3_8_1_bar CIM_cell
X2862 I382 O_3_8_2_2 WL_3_2 BL BLB W_3_8_2 W_3_8_2_bar CIM_cell
X2863 I382 O_3_8_2_3 WL_3_2 BL BLB W_3_8_3 W_3_8_3_bar CIM_cell
X2864 I382 O_3_8_2_4 WL_3_2 BL BLB W_3_8_4 W_3_8_4_bar CIM_cell
X2871 I383 O_3_8_3_1 WL_3_3 BL BLB W_3_8_1 W_3_8_1_bar CIM_cell
X2872 I383 O_3_8_3_2 WL_3_3 BL BLB W_3_8_2 W_3_8_2_bar CIM_cell
X2873 I383 O_3_8_3_3 WL_3_3 BL BLB W_3_8_3 W_3_8_3_bar CIM_cell
X2874 I383 O_3_8_3_4 WL_3_3 BL BLB W_3_8_4 W_3_8_4_bar CIM_cell
X2881 I384 O_3_8_4_1 WL_3_4 BL BLB W_3_8_1 W_3_8_1_bar CIM_cell
X2882 I384 O_3_8_4_2 WL_3_4 BL BLB W_3_8_2 W_3_8_2_bar CIM_cell
X2883 I384 O_3_8_4_3 WL_3_4 BL BLB W_3_8_3 W_3_8_3_bar CIM_cell
X2884 I384 O_3_8_4_4 WL_3_4 BL BLB W_3_8_4 W_3_8_4_bar CIM_cell
X2891 I391 O_3_9_1_1 WL_3_1 BL BLB W_3_9_1 W_3_9_1_bar CIM_cell
X2892 I391 O_3_9_1_2 WL_3_1 BL BLB W_3_9_2 W_3_9_2_bar CIM_cell
X2893 I391 O_3_9_1_3 WL_3_1 BL BLB W_3_9_3 W_3_9_3_bar CIM_cell
X2894 I391 O_3_9_1_4 WL_3_1 BL BLB W_3_9_4 W_3_9_4_bar CIM_cell
X2901 I392 O_3_9_2_1 WL_3_2 BL BLB W_3_9_1 W_3_9_1_bar CIM_cell
X2902 I392 O_3_9_2_2 WL_3_2 BL BLB W_3_9_2 W_3_9_2_bar CIM_cell
X2903 I392 O_3_9_2_3 WL_3_2 BL BLB W_3_9_3 W_3_9_3_bar CIM_cell
X2904 I392 O_3_9_2_4 WL_3_2 BL BLB W_3_9_4 W_3_9_4_bar CIM_cell
X2911 I393 O_3_9_3_1 WL_3_3 BL BLB W_3_9_1 W_3_9_1_bar CIM_cell
X2912 I393 O_3_9_3_2 WL_3_3 BL BLB W_3_9_2 W_3_9_2_bar CIM_cell
X2913 I393 O_3_9_3_3 WL_3_3 BL BLB W_3_9_3 W_3_9_3_bar CIM_cell
X2914 I393 O_3_9_3_4 WL_3_3 BL BLB W_3_9_4 W_3_9_4_bar CIM_cell
X2921 I394 O_3_9_4_1 WL_3_4 BL BLB W_3_9_1 W_3_9_1_bar CIM_cell
X2922 I394 O_3_9_4_2 WL_3_4 BL BLB W_3_9_2 W_3_9_2_bar CIM_cell
X2923 I394 O_3_9_4_3 WL_3_4 BL BLB W_3_9_3 W_3_9_3_bar CIM_cell
X2924 I394 O_3_9_4_4 WL_3_4 BL BLB W_3_9_4 W_3_9_4_bar CIM_cell
X2931 I3101 O_3_10_1_1 WL_3_1 BL BLB W_3_10_1 W_3_10_1_bar CIM_cell
X2932 I3101 O_3_10_1_2 WL_3_1 BL BLB W_3_10_2 W_3_10_2_bar CIM_cell
X2933 I3101 O_3_10_1_3 WL_3_1 BL BLB W_3_10_3 W_3_10_3_bar CIM_cell
X2934 I3101 O_3_10_1_4 WL_3_1 BL BLB W_3_10_4 W_3_10_4_bar CIM_cell
X2941 I3102 O_3_10_2_1 WL_3_2 BL BLB W_3_10_1 W_3_10_1_bar CIM_cell
X2942 I3102 O_3_10_2_2 WL_3_2 BL BLB W_3_10_2 W_3_10_2_bar CIM_cell
X2943 I3102 O_3_10_2_3 WL_3_2 BL BLB W_3_10_3 W_3_10_3_bar CIM_cell
X2944 I3102 O_3_10_2_4 WL_3_2 BL BLB W_3_10_4 W_3_10_4_bar CIM_cell
X2951 I3103 O_3_10_3_1 WL_3_3 BL BLB W_3_10_1 W_3_10_1_bar CIM_cell
X2952 I3103 O_3_10_3_2 WL_3_3 BL BLB W_3_10_2 W_3_10_2_bar CIM_cell
X2953 I3103 O_3_10_3_3 WL_3_3 BL BLB W_3_10_3 W_3_10_3_bar CIM_cell
X2954 I3103 O_3_10_3_4 WL_3_3 BL BLB W_3_10_4 W_3_10_4_bar CIM_cell
X2961 I3104 O_3_10_4_1 WL_3_4 BL BLB W_3_10_1 W_3_10_1_bar CIM_cell
X2962 I3104 O_3_10_4_2 WL_3_4 BL BLB W_3_10_2 W_3_10_2_bar CIM_cell
X2963 I3104 O_3_10_4_3 WL_3_4 BL BLB W_3_10_3 W_3_10_3_bar CIM_cell
X2964 I3104 O_3_10_4_4 WL_3_4 BL BLB W_3_10_4 W_3_10_4_bar CIM_cell
X2971 I3111 O_3_11_1_1 WL_3_1 BL BLB W_3_11_1 W_3_11_1_bar CIM_cell
X2972 I3111 O_3_11_1_2 WL_3_1 BL BLB W_3_11_2 W_3_11_2_bar CIM_cell
X2973 I3111 O_3_11_1_3 WL_3_1 BL BLB W_3_11_3 W_3_11_3_bar CIM_cell
X2974 I3111 O_3_11_1_4 WL_3_1 BL BLB W_3_11_4 W_3_11_4_bar CIM_cell
X2981 I3112 O_3_11_2_1 WL_3_2 BL BLB W_3_11_1 W_3_11_1_bar CIM_cell
X2982 I3112 O_3_11_2_2 WL_3_2 BL BLB W_3_11_2 W_3_11_2_bar CIM_cell
X2983 I3112 O_3_11_2_3 WL_3_2 BL BLB W_3_11_3 W_3_11_3_bar CIM_cell
X2984 I3112 O_3_11_2_4 WL_3_2 BL BLB W_3_11_4 W_3_11_4_bar CIM_cell
X2991 I3113 O_3_11_3_1 WL_3_3 BL BLB W_3_11_1 W_3_11_1_bar CIM_cell
X2992 I3113 O_3_11_3_2 WL_3_3 BL BLB W_3_11_2 W_3_11_2_bar CIM_cell
X2993 I3113 O_3_11_3_3 WL_3_3 BL BLB W_3_11_3 W_3_11_3_bar CIM_cell
X2994 I3113 O_3_11_3_4 WL_3_3 BL BLB W_3_11_4 W_3_11_4_bar CIM_cell
X3001 I3114 O_3_11_4_1 WL_3_4 BL BLB W_3_11_1 W_3_11_1_bar CIM_cell
X3002 I3114 O_3_11_4_2 WL_3_4 BL BLB W_3_11_2 W_3_11_2_bar CIM_cell
X3003 I3114 O_3_11_4_3 WL_3_4 BL BLB W_3_11_3 W_3_11_3_bar CIM_cell
X3004 I3114 O_3_11_4_4 WL_3_4 BL BLB W_3_11_4 W_3_11_4_bar CIM_cell
X3011 I3121 O_3_12_1_1 WL_3_1 BL BLB W_3_12_1 W_3_12_1_bar CIM_cell
X3012 I3121 O_3_12_1_2 WL_3_1 BL BLB W_3_12_2 W_3_12_2_bar CIM_cell
X3013 I3121 O_3_12_1_3 WL_3_1 BL BLB W_3_12_3 W_3_12_3_bar CIM_cell
X3014 I3121 O_3_12_1_4 WL_3_1 BL BLB W_3_12_4 W_3_12_4_bar CIM_cell
X3021 I3122 O_3_12_2_1 WL_3_2 BL BLB W_3_12_1 W_3_12_1_bar CIM_cell
X3022 I3122 O_3_12_2_2 WL_3_2 BL BLB W_3_12_2 W_3_12_2_bar CIM_cell
X3023 I3122 O_3_12_2_3 WL_3_2 BL BLB W_3_12_3 W_3_12_3_bar CIM_cell
X3024 I3122 O_3_12_2_4 WL_3_2 BL BLB W_3_12_4 W_3_12_4_bar CIM_cell
X3031 I3123 O_3_12_3_1 WL_3_3 BL BLB W_3_12_1 W_3_12_1_bar CIM_cell
X3032 I3123 O_3_12_3_2 WL_3_3 BL BLB W_3_12_2 W_3_12_2_bar CIM_cell
X3033 I3123 O_3_12_3_3 WL_3_3 BL BLB W_3_12_3 W_3_12_3_bar CIM_cell
X3034 I3123 O_3_12_3_4 WL_3_3 BL BLB W_3_12_4 W_3_12_4_bar CIM_cell
X3041 I3124 O_3_12_4_1 WL_3_4 BL BLB W_3_12_1 W_3_12_1_bar CIM_cell
X3042 I3124 O_3_12_4_2 WL_3_4 BL BLB W_3_12_2 W_3_12_2_bar CIM_cell
X3043 I3124 O_3_12_4_3 WL_3_4 BL BLB W_3_12_3 W_3_12_3_bar CIM_cell
X3044 I3124 O_3_12_4_4 WL_3_4 BL BLB W_3_12_4 W_3_12_4_bar CIM_cell
X3051 I3131 O_3_13_1_1 WL_3_1 BL BLB W_3_13_1 W_3_13_1_bar CIM_cell
X3052 I3131 O_3_13_1_2 WL_3_1 BL BLB W_3_13_2 W_3_13_2_bar CIM_cell
X3053 I3131 O_3_13_1_3 WL_3_1 BL BLB W_3_13_3 W_3_13_3_bar CIM_cell
X3054 I3131 O_3_13_1_4 WL_3_1 BL BLB W_3_13_4 W_3_13_4_bar CIM_cell
X3061 I3132 O_3_13_2_1 WL_3_2 BL BLB W_3_13_1 W_3_13_1_bar CIM_cell
X3062 I3132 O_3_13_2_2 WL_3_2 BL BLB W_3_13_2 W_3_13_2_bar CIM_cell
X3063 I3132 O_3_13_2_3 WL_3_2 BL BLB W_3_13_3 W_3_13_3_bar CIM_cell
X3064 I3132 O_3_13_2_4 WL_3_2 BL BLB W_3_13_4 W_3_13_4_bar CIM_cell
X3071 I3133 O_3_13_3_1 WL_3_3 BL BLB W_3_13_1 W_3_13_1_bar CIM_cell
X3072 I3133 O_3_13_3_2 WL_3_3 BL BLB W_3_13_2 W_3_13_2_bar CIM_cell
X3073 I3133 O_3_13_3_3 WL_3_3 BL BLB W_3_13_3 W_3_13_3_bar CIM_cell
X3074 I3133 O_3_13_3_4 WL_3_3 BL BLB W_3_13_4 W_3_13_4_bar CIM_cell
X3081 I3134 O_3_13_4_1 WL_3_4 BL BLB W_3_13_1 W_3_13_1_bar CIM_cell
X3082 I3134 O_3_13_4_2 WL_3_4 BL BLB W_3_13_2 W_3_13_2_bar CIM_cell
X3083 I3134 O_3_13_4_3 WL_3_4 BL BLB W_3_13_3 W_3_13_3_bar CIM_cell
X3084 I3134 O_3_13_4_4 WL_3_4 BL BLB W_3_13_4 W_3_13_4_bar CIM_cell
X3091 I3141 O_3_14_1_1 WL_3_1 BL BLB W_3_14_1 W_3_14_1_bar CIM_cell
X3092 I3141 O_3_14_1_2 WL_3_1 BL BLB W_3_14_2 W_3_14_2_bar CIM_cell
X3093 I3141 O_3_14_1_3 WL_3_1 BL BLB W_3_14_3 W_3_14_3_bar CIM_cell
X3094 I3141 O_3_14_1_4 WL_3_1 BL BLB W_3_14_4 W_3_14_4_bar CIM_cell
X3101 I3142 O_3_14_2_1 WL_3_2 BL BLB W_3_14_1 W_3_14_1_bar CIM_cell
X3102 I3142 O_3_14_2_2 WL_3_2 BL BLB W_3_14_2 W_3_14_2_bar CIM_cell
X3103 I3142 O_3_14_2_3 WL_3_2 BL BLB W_3_14_3 W_3_14_3_bar CIM_cell
X3104 I3142 O_3_14_2_4 WL_3_2 BL BLB W_3_14_4 W_3_14_4_bar CIM_cell
X3111 I3143 O_3_14_3_1 WL_3_3 BL BLB W_3_14_1 W_3_14_1_bar CIM_cell
X3112 I3143 O_3_14_3_2 WL_3_3 BL BLB W_3_14_2 W_3_14_2_bar CIM_cell
X3113 I3143 O_3_14_3_3 WL_3_3 BL BLB W_3_14_3 W_3_14_3_bar CIM_cell
X3114 I3143 O_3_14_3_4 WL_3_3 BL BLB W_3_14_4 W_3_14_4_bar CIM_cell
X3121 I3144 O_3_14_4_1 WL_3_4 BL BLB W_3_14_1 W_3_14_1_bar CIM_cell
X3122 I3144 O_3_14_4_2 WL_3_4 BL BLB W_3_14_2 W_3_14_2_bar CIM_cell
X3123 I3144 O_3_14_4_3 WL_3_4 BL BLB W_3_14_3 W_3_14_3_bar CIM_cell
X3124 I3144 O_3_14_4_4 WL_3_4 BL BLB W_3_14_4 W_3_14_4_bar CIM_cell
X3131 I3151 O_3_15_1_1 WL_3_1 BL BLB W_3_15_1 W_3_15_1_bar CIM_cell
X3132 I3151 O_3_15_1_2 WL_3_1 BL BLB W_3_15_2 W_3_15_2_bar CIM_cell
X3133 I3151 O_3_15_1_3 WL_3_1 BL BLB W_3_15_3 W_3_15_3_bar CIM_cell
X3134 I3151 O_3_15_1_4 WL_3_1 BL BLB W_3_15_4 W_3_15_4_bar CIM_cell
X3141 I3152 O_3_15_2_1 WL_3_2 BL BLB W_3_15_1 W_3_15_1_bar CIM_cell
X3142 I3152 O_3_15_2_2 WL_3_2 BL BLB W_3_15_2 W_3_15_2_bar CIM_cell
X3143 I3152 O_3_15_2_3 WL_3_2 BL BLB W_3_15_3 W_3_15_3_bar CIM_cell
X3144 I3152 O_3_15_2_4 WL_3_2 BL BLB W_3_15_4 W_3_15_4_bar CIM_cell
X3151 I3153 O_3_15_3_1 WL_3_3 BL BLB W_3_15_1 W_3_15_1_bar CIM_cell
X3152 I3153 O_3_15_3_2 WL_3_3 BL BLB W_3_15_2 W_3_15_2_bar CIM_cell
X3153 I3153 O_3_15_3_3 WL_3_3 BL BLB W_3_15_3 W_3_15_3_bar CIM_cell
X3154 I3153 O_3_15_3_4 WL_3_3 BL BLB W_3_15_4 W_3_15_4_bar CIM_cell
X3161 I3154 O_3_15_4_1 WL_3_4 BL BLB W_3_15_1 W_3_15_1_bar CIM_cell
X3162 I3154 O_3_15_4_2 WL_3_4 BL BLB W_3_15_2 W_3_15_2_bar CIM_cell
X3163 I3154 O_3_15_4_3 WL_3_4 BL BLB W_3_15_3 W_3_15_3_bar CIM_cell
X3164 I3154 O_3_15_4_4 WL_3_4 BL BLB W_3_15_4 W_3_15_4_bar CIM_cell
X3171 I3161 O_3_16_1_1 WL_3_1 BL BLB W_3_16_1 W_3_16_1_bar CIM_cell
X3172 I3161 O_3_16_1_2 WL_3_1 BL BLB W_3_16_2 W_3_16_2_bar CIM_cell
X3173 I3161 O_3_16_1_3 WL_3_1 BL BLB W_3_16_3 W_3_16_3_bar CIM_cell
X3174 I3161 O_3_16_1_4 WL_3_1 BL BLB W_3_16_4 W_3_16_4_bar CIM_cell
X3181 I3162 O_3_16_2_1 WL_3_2 BL BLB W_3_16_1 W_3_16_1_bar CIM_cell
X3182 I3162 O_3_16_2_2 WL_3_2 BL BLB W_3_16_2 W_3_16_2_bar CIM_cell
X3183 I3162 O_3_16_2_3 WL_3_2 BL BLB W_3_16_3 W_3_16_3_bar CIM_cell
X3184 I3162 O_3_16_2_4 WL_3_2 BL BLB W_3_16_4 W_3_16_4_bar CIM_cell
X3191 I3163 O_3_16_3_1 WL_3_3 BL BLB W_3_16_1 W_3_16_1_bar CIM_cell
X3192 I3163 O_3_16_3_2 WL_3_3 BL BLB W_3_16_2 W_3_16_2_bar CIM_cell
X3193 I3163 O_3_16_3_3 WL_3_3 BL BLB W_3_16_3 W_3_16_3_bar CIM_cell
X3194 I3163 O_3_16_3_4 WL_3_3 BL BLB W_3_16_4 W_3_16_4_bar CIM_cell
X3201 I3164 O_3_16_4_1 WL_3_4 BL BLB W_3_16_1 W_3_16_1_bar CIM_cell
X3202 I3164 O_3_16_4_2 WL_3_4 BL BLB W_3_16_2 W_3_16_2_bar CIM_cell
X3203 I3164 O_3_16_4_3 WL_3_4 BL BLB W_3_16_3 W_3_16_3_bar CIM_cell
X3204 I3164 O_3_16_4_4 WL_3_4 BL BLB W_3_16_4 W_3_16_4_bar CIM_cell
X3211 I3171 O_3_17_1_1 WL_3_1 BL BLB W_3_17_1 W_3_17_1_bar CIM_cell
X3212 I3171 O_3_17_1_2 WL_3_1 BL BLB W_3_17_2 W_3_17_2_bar CIM_cell
X3213 I3171 O_3_17_1_3 WL_3_1 BL BLB W_3_17_3 W_3_17_3_bar CIM_cell
X3214 I3171 O_3_17_1_4 WL_3_1 BL BLB W_3_17_4 W_3_17_4_bar CIM_cell
X3221 I3172 O_3_17_2_1 WL_3_2 BL BLB W_3_17_1 W_3_17_1_bar CIM_cell
X3222 I3172 O_3_17_2_2 WL_3_2 BL BLB W_3_17_2 W_3_17_2_bar CIM_cell
X3223 I3172 O_3_17_2_3 WL_3_2 BL BLB W_3_17_3 W_3_17_3_bar CIM_cell
X3224 I3172 O_3_17_2_4 WL_3_2 BL BLB W_3_17_4 W_3_17_4_bar CIM_cell
X3231 I3173 O_3_17_3_1 WL_3_3 BL BLB W_3_17_1 W_3_17_1_bar CIM_cell
X3232 I3173 O_3_17_3_2 WL_3_3 BL BLB W_3_17_2 W_3_17_2_bar CIM_cell
X3233 I3173 O_3_17_3_3 WL_3_3 BL BLB W_3_17_3 W_3_17_3_bar CIM_cell
X3234 I3173 O_3_17_3_4 WL_3_3 BL BLB W_3_17_4 W_3_17_4_bar CIM_cell
X3241 I3174 O_3_17_4_1 WL_3_4 BL BLB W_3_17_1 W_3_17_1_bar CIM_cell
X3242 I3174 O_3_17_4_2 WL_3_4 BL BLB W_3_17_2 W_3_17_2_bar CIM_cell
X3243 I3174 O_3_17_4_3 WL_3_4 BL BLB W_3_17_3 W_3_17_3_bar CIM_cell
X3244 I3174 O_3_17_4_4 WL_3_4 BL BLB W_3_17_4 W_3_17_4_bar CIM_cell
X3251 I3181 O_3_18_1_1 WL_3_1 BL BLB W_3_18_1 W_3_18_1_bar CIM_cell
X3252 I3181 O_3_18_1_2 WL_3_1 BL BLB W_3_18_2 W_3_18_2_bar CIM_cell
X3253 I3181 O_3_18_1_3 WL_3_1 BL BLB W_3_18_3 W_3_18_3_bar CIM_cell
X3254 I3181 O_3_18_1_4 WL_3_1 BL BLB W_3_18_4 W_3_18_4_bar CIM_cell
X3261 I3182 O_3_18_2_1 WL_3_2 BL BLB W_3_18_1 W_3_18_1_bar CIM_cell
X3262 I3182 O_3_18_2_2 WL_3_2 BL BLB W_3_18_2 W_3_18_2_bar CIM_cell
X3263 I3182 O_3_18_2_3 WL_3_2 BL BLB W_3_18_3 W_3_18_3_bar CIM_cell
X3264 I3182 O_3_18_2_4 WL_3_2 BL BLB W_3_18_4 W_3_18_4_bar CIM_cell
X3271 I3183 O_3_18_3_1 WL_3_3 BL BLB W_3_18_1 W_3_18_1_bar CIM_cell
X3272 I3183 O_3_18_3_2 WL_3_3 BL BLB W_3_18_2 W_3_18_2_bar CIM_cell
X3273 I3183 O_3_18_3_3 WL_3_3 BL BLB W_3_18_3 W_3_18_3_bar CIM_cell
X3274 I3183 O_3_18_3_4 WL_3_3 BL BLB W_3_18_4 W_3_18_4_bar CIM_cell
X3281 I3184 O_3_18_4_1 WL_3_4 BL BLB W_3_18_1 W_3_18_1_bar CIM_cell
X3282 I3184 O_3_18_4_2 WL_3_4 BL BLB W_3_18_2 W_3_18_2_bar CIM_cell
X3283 I3184 O_3_18_4_3 WL_3_4 BL BLB W_3_18_3 W_3_18_3_bar CIM_cell
X3284 I3184 O_3_18_4_4 WL_3_4 BL BLB W_3_18_4 W_3_18_4_bar CIM_cell
X3291 I3191 O_3_19_1_1 WL_3_1 BL BLB W_3_19_1 W_3_19_1_bar CIM_cell
X3292 I3191 O_3_19_1_2 WL_3_1 BL BLB W_3_19_2 W_3_19_2_bar CIM_cell
X3293 I3191 O_3_19_1_3 WL_3_1 BL BLB W_3_19_3 W_3_19_3_bar CIM_cell
X3294 I3191 O_3_19_1_4 WL_3_1 BL BLB W_3_19_4 W_3_19_4_bar CIM_cell
X3301 I3192 O_3_19_2_1 WL_3_2 BL BLB W_3_19_1 W_3_19_1_bar CIM_cell
X3302 I3192 O_3_19_2_2 WL_3_2 BL BLB W_3_19_2 W_3_19_2_bar CIM_cell
X3303 I3192 O_3_19_2_3 WL_3_2 BL BLB W_3_19_3 W_3_19_3_bar CIM_cell
X3304 I3192 O_3_19_2_4 WL_3_2 BL BLB W_3_19_4 W_3_19_4_bar CIM_cell
X3311 I3193 O_3_19_3_1 WL_3_3 BL BLB W_3_19_1 W_3_19_1_bar CIM_cell
X3312 I3193 O_3_19_3_2 WL_3_3 BL BLB W_3_19_2 W_3_19_2_bar CIM_cell
X3313 I3193 O_3_19_3_3 WL_3_3 BL BLB W_3_19_3 W_3_19_3_bar CIM_cell
X3314 I3193 O_3_19_3_4 WL_3_3 BL BLB W_3_19_4 W_3_19_4_bar CIM_cell
X3321 I3194 O_3_19_4_1 WL_3_4 BL BLB W_3_19_1 W_3_19_1_bar CIM_cell
X3322 I3194 O_3_19_4_2 WL_3_4 BL BLB W_3_19_2 W_3_19_2_bar CIM_cell
X3323 I3194 O_3_19_4_3 WL_3_4 BL BLB W_3_19_3 W_3_19_3_bar CIM_cell
X3324 I3194 O_3_19_4_4 WL_3_4 BL BLB W_3_19_4 W_3_19_4_bar CIM_cell
X3331 I3201 O_3_20_1_1 WL_3_1 BL BLB W_3_20_1 W_3_20_1_bar CIM_cell
X3332 I3201 O_3_20_1_2 WL_3_1 BL BLB W_3_20_2 W_3_20_2_bar CIM_cell
X3333 I3201 O_3_20_1_3 WL_3_1 BL BLB W_3_20_3 W_3_20_3_bar CIM_cell
X3334 I3201 O_3_20_1_4 WL_3_1 BL BLB W_3_20_4 W_3_20_4_bar CIM_cell
X3341 I3202 O_3_20_2_1 WL_3_2 BL BLB W_3_20_1 W_3_20_1_bar CIM_cell
X3342 I3202 O_3_20_2_2 WL_3_2 BL BLB W_3_20_2 W_3_20_2_bar CIM_cell
X3343 I3202 O_3_20_2_3 WL_3_2 BL BLB W_3_20_3 W_3_20_3_bar CIM_cell
X3344 I3202 O_3_20_2_4 WL_3_2 BL BLB W_3_20_4 W_3_20_4_bar CIM_cell
X3351 I3203 O_3_20_3_1 WL_3_3 BL BLB W_3_20_1 W_3_20_1_bar CIM_cell
X3352 I3203 O_3_20_3_2 WL_3_3 BL BLB W_3_20_2 W_3_20_2_bar CIM_cell
X3353 I3203 O_3_20_3_3 WL_3_3 BL BLB W_3_20_3 W_3_20_3_bar CIM_cell
X3354 I3203 O_3_20_3_4 WL_3_3 BL BLB W_3_20_4 W_3_20_4_bar CIM_cell
X3361 I3204 O_3_20_4_1 WL_3_4 BL BLB W_3_20_1 W_3_20_1_bar CIM_cell
X3362 I3204 O_3_20_4_2 WL_3_4 BL BLB W_3_20_2 W_3_20_2_bar CIM_cell
X3363 I3204 O_3_20_4_3 WL_3_4 BL BLB W_3_20_3 W_3_20_3_bar CIM_cell
X3364 I3204 O_3_20_4_4 WL_3_4 BL BLB W_3_20_4 W_3_20_4_bar CIM_cell
X3371 I3211 O_3_21_1_1 WL_3_1 BL BLB W_3_21_1 W_3_21_1_bar CIM_cell
X3372 I3211 O_3_21_1_2 WL_3_1 BL BLB W_3_21_2 W_3_21_2_bar CIM_cell
X3373 I3211 O_3_21_1_3 WL_3_1 BL BLB W_3_21_3 W_3_21_3_bar CIM_cell
X3374 I3211 O_3_21_1_4 WL_3_1 BL BLB W_3_21_4 W_3_21_4_bar CIM_cell
X3381 I3212 O_3_21_2_1 WL_3_2 BL BLB W_3_21_1 W_3_21_1_bar CIM_cell
X3382 I3212 O_3_21_2_2 WL_3_2 BL BLB W_3_21_2 W_3_21_2_bar CIM_cell
X3383 I3212 O_3_21_2_3 WL_3_2 BL BLB W_3_21_3 W_3_21_3_bar CIM_cell
X3384 I3212 O_3_21_2_4 WL_3_2 BL BLB W_3_21_4 W_3_21_4_bar CIM_cell
X3391 I3213 O_3_21_3_1 WL_3_3 BL BLB W_3_21_1 W_3_21_1_bar CIM_cell
X3392 I3213 O_3_21_3_2 WL_3_3 BL BLB W_3_21_2 W_3_21_2_bar CIM_cell
X3393 I3213 O_3_21_3_3 WL_3_3 BL BLB W_3_21_3 W_3_21_3_bar CIM_cell
X3394 I3213 O_3_21_3_4 WL_3_3 BL BLB W_3_21_4 W_3_21_4_bar CIM_cell
X3401 I3214 O_3_21_4_1 WL_3_4 BL BLB W_3_21_1 W_3_21_1_bar CIM_cell
X3402 I3214 O_3_21_4_2 WL_3_4 BL BLB W_3_21_2 W_3_21_2_bar CIM_cell
X3403 I3214 O_3_21_4_3 WL_3_4 BL BLB W_3_21_3 W_3_21_3_bar CIM_cell
X3404 I3214 O_3_21_4_4 WL_3_4 BL BLB W_3_21_4 W_3_21_4_bar CIM_cell
X3411 I3221 O_3_22_1_1 WL_3_1 BL BLB W_3_22_1 W_3_22_1_bar CIM_cell
X3412 I3221 O_3_22_1_2 WL_3_1 BL BLB W_3_22_2 W_3_22_2_bar CIM_cell
X3413 I3221 O_3_22_1_3 WL_3_1 BL BLB W_3_22_3 W_3_22_3_bar CIM_cell
X3414 I3221 O_3_22_1_4 WL_3_1 BL BLB W_3_22_4 W_3_22_4_bar CIM_cell
X3421 I3222 O_3_22_2_1 WL_3_2 BL BLB W_3_22_1 W_3_22_1_bar CIM_cell
X3422 I3222 O_3_22_2_2 WL_3_2 BL BLB W_3_22_2 W_3_22_2_bar CIM_cell
X3423 I3222 O_3_22_2_3 WL_3_2 BL BLB W_3_22_3 W_3_22_3_bar CIM_cell
X3424 I3222 O_3_22_2_4 WL_3_2 BL BLB W_3_22_4 W_3_22_4_bar CIM_cell
X3431 I3223 O_3_22_3_1 WL_3_3 BL BLB W_3_22_1 W_3_22_1_bar CIM_cell
X3432 I3223 O_3_22_3_2 WL_3_3 BL BLB W_3_22_2 W_3_22_2_bar CIM_cell
X3433 I3223 O_3_22_3_3 WL_3_3 BL BLB W_3_22_3 W_3_22_3_bar CIM_cell
X3434 I3223 O_3_22_3_4 WL_3_3 BL BLB W_3_22_4 W_3_22_4_bar CIM_cell
X3441 I3224 O_3_22_4_1 WL_3_4 BL BLB W_3_22_1 W_3_22_1_bar CIM_cell
X3442 I3224 O_3_22_4_2 WL_3_4 BL BLB W_3_22_2 W_3_22_2_bar CIM_cell
X3443 I3224 O_3_22_4_3 WL_3_4 BL BLB W_3_22_3 W_3_22_3_bar CIM_cell
X3444 I3224 O_3_22_4_4 WL_3_4 BL BLB W_3_22_4 W_3_22_4_bar CIM_cell
X3451 I3231 O_3_23_1_1 WL_3_1 BL BLB W_3_23_1 W_3_23_1_bar CIM_cell
X3452 I3231 O_3_23_1_2 WL_3_1 BL BLB W_3_23_2 W_3_23_2_bar CIM_cell
X3453 I3231 O_3_23_1_3 WL_3_1 BL BLB W_3_23_3 W_3_23_3_bar CIM_cell
X3454 I3231 O_3_23_1_4 WL_3_1 BL BLB W_3_23_4 W_3_23_4_bar CIM_cell
X3461 I3232 O_3_23_2_1 WL_3_2 BL BLB W_3_23_1 W_3_23_1_bar CIM_cell
X3462 I3232 O_3_23_2_2 WL_3_2 BL BLB W_3_23_2 W_3_23_2_bar CIM_cell
X3463 I3232 O_3_23_2_3 WL_3_2 BL BLB W_3_23_3 W_3_23_3_bar CIM_cell
X3464 I3232 O_3_23_2_4 WL_3_2 BL BLB W_3_23_4 W_3_23_4_bar CIM_cell
X3471 I3233 O_3_23_3_1 WL_3_3 BL BLB W_3_23_1 W_3_23_1_bar CIM_cell
X3472 I3233 O_3_23_3_2 WL_3_3 BL BLB W_3_23_2 W_3_23_2_bar CIM_cell
X3473 I3233 O_3_23_3_3 WL_3_3 BL BLB W_3_23_3 W_3_23_3_bar CIM_cell
X3474 I3233 O_3_23_3_4 WL_3_3 BL BLB W_3_23_4 W_3_23_4_bar CIM_cell
X3481 I3234 O_3_23_4_1 WL_3_4 BL BLB W_3_23_1 W_3_23_1_bar CIM_cell
X3482 I3234 O_3_23_4_2 WL_3_4 BL BLB W_3_23_2 W_3_23_2_bar CIM_cell
X3483 I3234 O_3_23_4_3 WL_3_4 BL BLB W_3_23_3 W_3_23_3_bar CIM_cell
X3484 I3234 O_3_23_4_4 WL_3_4 BL BLB W_3_23_4 W_3_23_4_bar CIM_cell
X3491 I3241 O_3_24_1_1 WL_3_1 BL BLB W_3_24_1 W_3_24_1_bar CIM_cell
X3492 I3241 O_3_24_1_2 WL_3_1 BL BLB W_3_24_2 W_3_24_2_bar CIM_cell
X3493 I3241 O_3_24_1_3 WL_3_1 BL BLB W_3_24_3 W_3_24_3_bar CIM_cell
X3494 I3241 O_3_24_1_4 WL_3_1 BL BLB W_3_24_4 W_3_24_4_bar CIM_cell
X3501 I3242 O_3_24_2_1 WL_3_2 BL BLB W_3_24_1 W_3_24_1_bar CIM_cell
X3502 I3242 O_3_24_2_2 WL_3_2 BL BLB W_3_24_2 W_3_24_2_bar CIM_cell
X3503 I3242 O_3_24_2_3 WL_3_2 BL BLB W_3_24_3 W_3_24_3_bar CIM_cell
X3504 I3242 O_3_24_2_4 WL_3_2 BL BLB W_3_24_4 W_3_24_4_bar CIM_cell
X3511 I3243 O_3_24_3_1 WL_3_3 BL BLB W_3_24_1 W_3_24_1_bar CIM_cell
X3512 I3243 O_3_24_3_2 WL_3_3 BL BLB W_3_24_2 W_3_24_2_bar CIM_cell
X3513 I3243 O_3_24_3_3 WL_3_3 BL BLB W_3_24_3 W_3_24_3_bar CIM_cell
X3514 I3243 O_3_24_3_4 WL_3_3 BL BLB W_3_24_4 W_3_24_4_bar CIM_cell
X3521 I3244 O_3_24_4_1 WL_3_4 BL BLB W_3_24_1 W_3_24_1_bar CIM_cell
X3522 I3244 O_3_24_4_2 WL_3_4 BL BLB W_3_24_2 W_3_24_2_bar CIM_cell
X3523 I3244 O_3_24_4_3 WL_3_4 BL BLB W_3_24_3 W_3_24_3_bar CIM_cell
X3524 I3244 O_3_24_4_4 WL_3_4 BL BLB W_3_24_4 W_3_24_4_bar CIM_cell
X3531 I3251 O_3_25_1_1 WL_3_1 BL BLB W_3_25_1 W_3_25_1_bar CIM_cell
X3532 I3251 O_3_25_1_2 WL_3_1 BL BLB W_3_25_2 W_3_25_2_bar CIM_cell
X3533 I3251 O_3_25_1_3 WL_3_1 BL BLB W_3_25_3 W_3_25_3_bar CIM_cell
X3534 I3251 O_3_25_1_4 WL_3_1 BL BLB W_3_25_4 W_3_25_4_bar CIM_cell
X3541 I3252 O_3_25_2_1 WL_3_2 BL BLB W_3_25_1 W_3_25_1_bar CIM_cell
X3542 I3252 O_3_25_2_2 WL_3_2 BL BLB W_3_25_2 W_3_25_2_bar CIM_cell
X3543 I3252 O_3_25_2_3 WL_3_2 BL BLB W_3_25_3 W_3_25_3_bar CIM_cell
X3544 I3252 O_3_25_2_4 WL_3_2 BL BLB W_3_25_4 W_3_25_4_bar CIM_cell
X3551 I3253 O_3_25_3_1 WL_3_3 BL BLB W_3_25_1 W_3_25_1_bar CIM_cell
X3552 I3253 O_3_25_3_2 WL_3_3 BL BLB W_3_25_2 W_3_25_2_bar CIM_cell
X3553 I3253 O_3_25_3_3 WL_3_3 BL BLB W_3_25_3 W_3_25_3_bar CIM_cell
X3554 I3253 O_3_25_3_4 WL_3_3 BL BLB W_3_25_4 W_3_25_4_bar CIM_cell
X3561 I3254 O_3_25_4_1 WL_3_4 BL BLB W_3_25_1 W_3_25_1_bar CIM_cell
X3562 I3254 O_3_25_4_2 WL_3_4 BL BLB W_3_25_2 W_3_25_2_bar CIM_cell
X3563 I3254 O_3_25_4_3 WL_3_4 BL BLB W_3_25_3 W_3_25_3_bar CIM_cell
X3564 I3254 O_3_25_4_4 WL_3_4 BL BLB W_3_25_4 W_3_25_4_bar CIM_cell
X3571 I3261 O_3_26_1_1 WL_3_1 BL BLB W_3_26_1 W_3_26_1_bar CIM_cell
X3572 I3261 O_3_26_1_2 WL_3_1 BL BLB W_3_26_2 W_3_26_2_bar CIM_cell
X3573 I3261 O_3_26_1_3 WL_3_1 BL BLB W_3_26_3 W_3_26_3_bar CIM_cell
X3574 I3261 O_3_26_1_4 WL_3_1 BL BLB W_3_26_4 W_3_26_4_bar CIM_cell
X3581 I3262 O_3_26_2_1 WL_3_2 BL BLB W_3_26_1 W_3_26_1_bar CIM_cell
X3582 I3262 O_3_26_2_2 WL_3_2 BL BLB W_3_26_2 W_3_26_2_bar CIM_cell
X3583 I3262 O_3_26_2_3 WL_3_2 BL BLB W_3_26_3 W_3_26_3_bar CIM_cell
X3584 I3262 O_3_26_2_4 WL_3_2 BL BLB W_3_26_4 W_3_26_4_bar CIM_cell
X3591 I3263 O_3_26_3_1 WL_3_3 BL BLB W_3_26_1 W_3_26_1_bar CIM_cell
X3592 I3263 O_3_26_3_2 WL_3_3 BL BLB W_3_26_2 W_3_26_2_bar CIM_cell
X3593 I3263 O_3_26_3_3 WL_3_3 BL BLB W_3_26_3 W_3_26_3_bar CIM_cell
X3594 I3263 O_3_26_3_4 WL_3_3 BL BLB W_3_26_4 W_3_26_4_bar CIM_cell
X3601 I3264 O_3_26_4_1 WL_3_4 BL BLB W_3_26_1 W_3_26_1_bar CIM_cell
X3602 I3264 O_3_26_4_2 WL_3_4 BL BLB W_3_26_2 W_3_26_2_bar CIM_cell
X3603 I3264 O_3_26_4_3 WL_3_4 BL BLB W_3_26_3 W_3_26_3_bar CIM_cell
X3604 I3264 O_3_26_4_4 WL_3_4 BL BLB W_3_26_4 W_3_26_4_bar CIM_cell
X3611 I3271 O_3_27_1_1 WL_3_1 BL BLB W_3_27_1 W_3_27_1_bar CIM_cell
X3612 I3271 O_3_27_1_2 WL_3_1 BL BLB W_3_27_2 W_3_27_2_bar CIM_cell
X3613 I3271 O_3_27_1_3 WL_3_1 BL BLB W_3_27_3 W_3_27_3_bar CIM_cell
X3614 I3271 O_3_27_1_4 WL_3_1 BL BLB W_3_27_4 W_3_27_4_bar CIM_cell
X3621 I3272 O_3_27_2_1 WL_3_2 BL BLB W_3_27_1 W_3_27_1_bar CIM_cell
X3622 I3272 O_3_27_2_2 WL_3_2 BL BLB W_3_27_2 W_3_27_2_bar CIM_cell
X3623 I3272 O_3_27_2_3 WL_3_2 BL BLB W_3_27_3 W_3_27_3_bar CIM_cell
X3624 I3272 O_3_27_2_4 WL_3_2 BL BLB W_3_27_4 W_3_27_4_bar CIM_cell
X3631 I3273 O_3_27_3_1 WL_3_3 BL BLB W_3_27_1 W_3_27_1_bar CIM_cell
X3632 I3273 O_3_27_3_2 WL_3_3 BL BLB W_3_27_2 W_3_27_2_bar CIM_cell
X3633 I3273 O_3_27_3_3 WL_3_3 BL BLB W_3_27_3 W_3_27_3_bar CIM_cell
X3634 I3273 O_3_27_3_4 WL_3_3 BL BLB W_3_27_4 W_3_27_4_bar CIM_cell
X3641 I3274 O_3_27_4_1 WL_3_4 BL BLB W_3_27_1 W_3_27_1_bar CIM_cell
X3642 I3274 O_3_27_4_2 WL_3_4 BL BLB W_3_27_2 W_3_27_2_bar CIM_cell
X3643 I3274 O_3_27_4_3 WL_3_4 BL BLB W_3_27_3 W_3_27_3_bar CIM_cell
X3644 I3274 O_3_27_4_4 WL_3_4 BL BLB W_3_27_4 W_3_27_4_bar CIM_cell
X3651 I3281 O_3_28_1_1 WL_3_1 BL BLB W_3_28_1 W_3_28_1_bar CIM_cell
X3652 I3281 O_3_28_1_2 WL_3_1 BL BLB W_3_28_2 W_3_28_2_bar CIM_cell
X3653 I3281 O_3_28_1_3 WL_3_1 BL BLB W_3_28_3 W_3_28_3_bar CIM_cell
X3654 I3281 O_3_28_1_4 WL_3_1 BL BLB W_3_28_4 W_3_28_4_bar CIM_cell
X3661 I3282 O_3_28_2_1 WL_3_2 BL BLB W_3_28_1 W_3_28_1_bar CIM_cell
X3662 I3282 O_3_28_2_2 WL_3_2 BL BLB W_3_28_2 W_3_28_2_bar CIM_cell
X3663 I3282 O_3_28_2_3 WL_3_2 BL BLB W_3_28_3 W_3_28_3_bar CIM_cell
X3664 I3282 O_3_28_2_4 WL_3_2 BL BLB W_3_28_4 W_3_28_4_bar CIM_cell
X3671 I3283 O_3_28_3_1 WL_3_3 BL BLB W_3_28_1 W_3_28_1_bar CIM_cell
X3672 I3283 O_3_28_3_2 WL_3_3 BL BLB W_3_28_2 W_3_28_2_bar CIM_cell
X3673 I3283 O_3_28_3_3 WL_3_3 BL BLB W_3_28_3 W_3_28_3_bar CIM_cell
X3674 I3283 O_3_28_3_4 WL_3_3 BL BLB W_3_28_4 W_3_28_4_bar CIM_cell
X3681 I3284 O_3_28_4_1 WL_3_4 BL BLB W_3_28_1 W_3_28_1_bar CIM_cell
X3682 I3284 O_3_28_4_2 WL_3_4 BL BLB W_3_28_2 W_3_28_2_bar CIM_cell
X3683 I3284 O_3_28_4_3 WL_3_4 BL BLB W_3_28_3 W_3_28_3_bar CIM_cell
X3684 I3284 O_3_28_4_4 WL_3_4 BL BLB W_3_28_4 W_3_28_4_bar CIM_cell
X3691 I3291 O_3_29_1_1 WL_3_1 BL BLB W_3_29_1 W_3_29_1_bar CIM_cell
X3692 I3291 O_3_29_1_2 WL_3_1 BL BLB W_3_29_2 W_3_29_2_bar CIM_cell
X3693 I3291 O_3_29_1_3 WL_3_1 BL BLB W_3_29_3 W_3_29_3_bar CIM_cell
X3694 I3291 O_3_29_1_4 WL_3_1 BL BLB W_3_29_4 W_3_29_4_bar CIM_cell
X3701 I3292 O_3_29_2_1 WL_3_2 BL BLB W_3_29_1 W_3_29_1_bar CIM_cell
X3702 I3292 O_3_29_2_2 WL_3_2 BL BLB W_3_29_2 W_3_29_2_bar CIM_cell
X3703 I3292 O_3_29_2_3 WL_3_2 BL BLB W_3_29_3 W_3_29_3_bar CIM_cell
X3704 I3292 O_3_29_2_4 WL_3_2 BL BLB W_3_29_4 W_3_29_4_bar CIM_cell
X3711 I3293 O_3_29_3_1 WL_3_3 BL BLB W_3_29_1 W_3_29_1_bar CIM_cell
X3712 I3293 O_3_29_3_2 WL_3_3 BL BLB W_3_29_2 W_3_29_2_bar CIM_cell
X3713 I3293 O_3_29_3_3 WL_3_3 BL BLB W_3_29_3 W_3_29_3_bar CIM_cell
X3714 I3293 O_3_29_3_4 WL_3_3 BL BLB W_3_29_4 W_3_29_4_bar CIM_cell
X3721 I3294 O_3_29_4_1 WL_3_4 BL BLB W_3_29_1 W_3_29_1_bar CIM_cell
X3722 I3294 O_3_29_4_2 WL_3_4 BL BLB W_3_29_2 W_3_29_2_bar CIM_cell
X3723 I3294 O_3_29_4_3 WL_3_4 BL BLB W_3_29_3 W_3_29_3_bar CIM_cell
X3724 I3294 O_3_29_4_4 WL_3_4 BL BLB W_3_29_4 W_3_29_4_bar CIM_cell
X3731 I3301 O_3_30_1_1 WL_3_1 BL BLB W_3_30_1 W_3_30_1_bar CIM_cell
X3732 I3301 O_3_30_1_2 WL_3_1 BL BLB W_3_30_2 W_3_30_2_bar CIM_cell
X3733 I3301 O_3_30_1_3 WL_3_1 BL BLB W_3_30_3 W_3_30_3_bar CIM_cell
X3734 I3301 O_3_30_1_4 WL_3_1 BL BLB W_3_30_4 W_3_30_4_bar CIM_cell
X3741 I3302 O_3_30_2_1 WL_3_2 BL BLB W_3_30_1 W_3_30_1_bar CIM_cell
X3742 I3302 O_3_30_2_2 WL_3_2 BL BLB W_3_30_2 W_3_30_2_bar CIM_cell
X3743 I3302 O_3_30_2_3 WL_3_2 BL BLB W_3_30_3 W_3_30_3_bar CIM_cell
X3744 I3302 O_3_30_2_4 WL_3_2 BL BLB W_3_30_4 W_3_30_4_bar CIM_cell
X3751 I3303 O_3_30_3_1 WL_3_3 BL BLB W_3_30_1 W_3_30_1_bar CIM_cell
X3752 I3303 O_3_30_3_2 WL_3_3 BL BLB W_3_30_2 W_3_30_2_bar CIM_cell
X3753 I3303 O_3_30_3_3 WL_3_3 BL BLB W_3_30_3 W_3_30_3_bar CIM_cell
X3754 I3303 O_3_30_3_4 WL_3_3 BL BLB W_3_30_4 W_3_30_4_bar CIM_cell
X3761 I3304 O_3_30_4_1 WL_3_4 BL BLB W_3_30_1 W_3_30_1_bar CIM_cell
X3762 I3304 O_3_30_4_2 WL_3_4 BL BLB W_3_30_2 W_3_30_2_bar CIM_cell
X3763 I3304 O_3_30_4_3 WL_3_4 BL BLB W_3_30_3 W_3_30_3_bar CIM_cell
X3764 I3304 O_3_30_4_4 WL_3_4 BL BLB W_3_30_4 W_3_30_4_bar CIM_cell
X3771 I3311 O_3_31_1_1 WL_3_1 BL BLB W_3_31_1 W_3_31_1_bar CIM_cell
X3772 I3311 O_3_31_1_2 WL_3_1 BL BLB W_3_31_2 W_3_31_2_bar CIM_cell
X3773 I3311 O_3_31_1_3 WL_3_1 BL BLB W_3_31_3 W_3_31_3_bar CIM_cell
X3774 I3311 O_3_31_1_4 WL_3_1 BL BLB W_3_31_4 W_3_31_4_bar CIM_cell
X3781 I3312 O_3_31_2_1 WL_3_2 BL BLB W_3_31_1 W_3_31_1_bar CIM_cell
X3782 I3312 O_3_31_2_2 WL_3_2 BL BLB W_3_31_2 W_3_31_2_bar CIM_cell
X3783 I3312 O_3_31_2_3 WL_3_2 BL BLB W_3_31_3 W_3_31_3_bar CIM_cell
X3784 I3312 O_3_31_2_4 WL_3_2 BL BLB W_3_31_4 W_3_31_4_bar CIM_cell
X3791 I3313 O_3_31_3_1 WL_3_3 BL BLB W_3_31_1 W_3_31_1_bar CIM_cell
X3792 I3313 O_3_31_3_2 WL_3_3 BL BLB W_3_31_2 W_3_31_2_bar CIM_cell
X3793 I3313 O_3_31_3_3 WL_3_3 BL BLB W_3_31_3 W_3_31_3_bar CIM_cell
X3794 I3313 O_3_31_3_4 WL_3_3 BL BLB W_3_31_4 W_3_31_4_bar CIM_cell
X3801 I3314 O_3_31_4_1 WL_3_4 BL BLB W_3_31_1 W_3_31_1_bar CIM_cell
X3802 I3314 O_3_31_4_2 WL_3_4 BL BLB W_3_31_2 W_3_31_2_bar CIM_cell
X3803 I3314 O_3_31_4_3 WL_3_4 BL BLB W_3_31_3 W_3_31_3_bar CIM_cell
X3804 I3314 O_3_31_4_4 WL_3_4 BL BLB W_3_31_4 W_3_31_4_bar CIM_cell
X3811 I3321 O_3_32_1_1 WL_3_1 BL BLB W_3_32_1 W_3_32_1_bar CIM_cell
X3812 I3321 O_3_32_1_2 WL_3_1 BL BLB W_3_32_2 W_3_32_2_bar CIM_cell
X3813 I3321 O_3_32_1_3 WL_3_1 BL BLB W_3_32_3 W_3_32_3_bar CIM_cell
X3814 I3321 O_3_32_1_4 WL_3_1 BL BLB W_3_32_4 W_3_32_4_bar CIM_cell
X3821 I3322 O_3_32_2_1 WL_3_2 BL BLB W_3_32_1 W_3_32_1_bar CIM_cell
X3822 I3322 O_3_32_2_2 WL_3_2 BL BLB W_3_32_2 W_3_32_2_bar CIM_cell
X3823 I3322 O_3_32_2_3 WL_3_2 BL BLB W_3_32_3 W_3_32_3_bar CIM_cell
X3824 I3322 O_3_32_2_4 WL_3_2 BL BLB W_3_32_4 W_3_32_4_bar CIM_cell
X3831 I3323 O_3_32_3_1 WL_3_3 BL BLB W_3_32_1 W_3_32_1_bar CIM_cell
X3832 I3323 O_3_32_3_2 WL_3_3 BL BLB W_3_32_2 W_3_32_2_bar CIM_cell
X3833 I3323 O_3_32_3_3 WL_3_3 BL BLB W_3_32_3 W_3_32_3_bar CIM_cell
X3834 I3323 O_3_32_3_4 WL_3_3 BL BLB W_3_32_4 W_3_32_4_bar CIM_cell
X3841 I3324 O_3_32_4_1 WL_3_4 BL BLB W_3_32_1 W_3_32_1_bar CIM_cell
X3842 I3324 O_3_32_4_2 WL_3_4 BL BLB W_3_32_2 W_3_32_2_bar CIM_cell
X3843 I3324 O_3_32_4_3 WL_3_4 BL BLB W_3_32_3 W_3_32_3_bar CIM_cell
X3844 I3324 O_3_32_4_4 WL_3_4 BL BLB W_3_32_4 W_3_32_4_bar CIM_cell
X3851 I411 O_4_1_1_1 WL_4_1 BL BLB W_4_1_1 W_4_1_1_bar CIM_cell
X3852 I411 O_4_1_1_2 WL_4_1 BL BLB W_4_1_2 W_4_1_2_bar CIM_cell
X3853 I411 O_4_1_1_3 WL_4_1 BL BLB W_4_1_3 W_4_1_3_bar CIM_cell
X3854 I411 O_4_1_1_4 WL_4_1 BL BLB W_4_1_4 W_4_1_4_bar CIM_cell
X3861 I412 O_4_1_2_1 WL_4_2 BL BLB W_4_1_1 W_4_1_1_bar CIM_cell
X3862 I412 O_4_1_2_2 WL_4_2 BL BLB W_4_1_2 W_4_1_2_bar CIM_cell
X3863 I412 O_4_1_2_3 WL_4_2 BL BLB W_4_1_3 W_4_1_3_bar CIM_cell
X3864 I412 O_4_1_2_4 WL_4_2 BL BLB W_4_1_4 W_4_1_4_bar CIM_cell
X3871 I413 O_4_1_3_1 WL_4_3 BL BLB W_4_1_1 W_4_1_1_bar CIM_cell
X3872 I413 O_4_1_3_2 WL_4_3 BL BLB W_4_1_2 W_4_1_2_bar CIM_cell
X3873 I413 O_4_1_3_3 WL_4_3 BL BLB W_4_1_3 W_4_1_3_bar CIM_cell
X3874 I413 O_4_1_3_4 WL_4_3 BL BLB W_4_1_4 W_4_1_4_bar CIM_cell
X3881 I414 O_4_1_4_1 WL_4_4 BL BLB W_4_1_1 W_4_1_1_bar CIM_cell
X3882 I414 O_4_1_4_2 WL_4_4 BL BLB W_4_1_2 W_4_1_2_bar CIM_cell
X3883 I414 O_4_1_4_3 WL_4_4 BL BLB W_4_1_3 W_4_1_3_bar CIM_cell
X3884 I414 O_4_1_4_4 WL_4_4 BL BLB W_4_1_4 W_4_1_4_bar CIM_cell
X3891 I421 O_4_2_1_1 WL_4_1 BL BLB W_4_2_1 W_4_2_1_bar CIM_cell
X3892 I421 O_4_2_1_2 WL_4_1 BL BLB W_4_2_2 W_4_2_2_bar CIM_cell
X3893 I421 O_4_2_1_3 WL_4_1 BL BLB W_4_2_3 W_4_2_3_bar CIM_cell
X3894 I421 O_4_2_1_4 WL_4_1 BL BLB W_4_2_4 W_4_2_4_bar CIM_cell
X3901 I422 O_4_2_2_1 WL_4_2 BL BLB W_4_2_1 W_4_2_1_bar CIM_cell
X3902 I422 O_4_2_2_2 WL_4_2 BL BLB W_4_2_2 W_4_2_2_bar CIM_cell
X3903 I422 O_4_2_2_3 WL_4_2 BL BLB W_4_2_3 W_4_2_3_bar CIM_cell
X3904 I422 O_4_2_2_4 WL_4_2 BL BLB W_4_2_4 W_4_2_4_bar CIM_cell
X3911 I423 O_4_2_3_1 WL_4_3 BL BLB W_4_2_1 W_4_2_1_bar CIM_cell
X3912 I423 O_4_2_3_2 WL_4_3 BL BLB W_4_2_2 W_4_2_2_bar CIM_cell
X3913 I423 O_4_2_3_3 WL_4_3 BL BLB W_4_2_3 W_4_2_3_bar CIM_cell
X3914 I423 O_4_2_3_4 WL_4_3 BL BLB W_4_2_4 W_4_2_4_bar CIM_cell
X3921 I424 O_4_2_4_1 WL_4_4 BL BLB W_4_2_1 W_4_2_1_bar CIM_cell
X3922 I424 O_4_2_4_2 WL_4_4 BL BLB W_4_2_2 W_4_2_2_bar CIM_cell
X3923 I424 O_4_2_4_3 WL_4_4 BL BLB W_4_2_3 W_4_2_3_bar CIM_cell
X3924 I424 O_4_2_4_4 WL_4_4 BL BLB W_4_2_4 W_4_2_4_bar CIM_cell
X3931 I431 O_4_3_1_1 WL_4_1 BL BLB W_4_3_1 W_4_3_1_bar CIM_cell
X3932 I431 O_4_3_1_2 WL_4_1 BL BLB W_4_3_2 W_4_3_2_bar CIM_cell
X3933 I431 O_4_3_1_3 WL_4_1 BL BLB W_4_3_3 W_4_3_3_bar CIM_cell
X3934 I431 O_4_3_1_4 WL_4_1 BL BLB W_4_3_4 W_4_3_4_bar CIM_cell
X3941 I432 O_4_3_2_1 WL_4_2 BL BLB W_4_3_1 W_4_3_1_bar CIM_cell
X3942 I432 O_4_3_2_2 WL_4_2 BL BLB W_4_3_2 W_4_3_2_bar CIM_cell
X3943 I432 O_4_3_2_3 WL_4_2 BL BLB W_4_3_3 W_4_3_3_bar CIM_cell
X3944 I432 O_4_3_2_4 WL_4_2 BL BLB W_4_3_4 W_4_3_4_bar CIM_cell
X3951 I433 O_4_3_3_1 WL_4_3 BL BLB W_4_3_1 W_4_3_1_bar CIM_cell
X3952 I433 O_4_3_3_2 WL_4_3 BL BLB W_4_3_2 W_4_3_2_bar CIM_cell
X3953 I433 O_4_3_3_3 WL_4_3 BL BLB W_4_3_3 W_4_3_3_bar CIM_cell
X3954 I433 O_4_3_3_4 WL_4_3 BL BLB W_4_3_4 W_4_3_4_bar CIM_cell
X3961 I434 O_4_3_4_1 WL_4_4 BL BLB W_4_3_1 W_4_3_1_bar CIM_cell
X3962 I434 O_4_3_4_2 WL_4_4 BL BLB W_4_3_2 W_4_3_2_bar CIM_cell
X3963 I434 O_4_3_4_3 WL_4_4 BL BLB W_4_3_3 W_4_3_3_bar CIM_cell
X3964 I434 O_4_3_4_4 WL_4_4 BL BLB W_4_3_4 W_4_3_4_bar CIM_cell
X3971 I441 O_4_4_1_1 WL_4_1 BL BLB W_4_4_1 W_4_4_1_bar CIM_cell
X3972 I441 O_4_4_1_2 WL_4_1 BL BLB W_4_4_2 W_4_4_2_bar CIM_cell
X3973 I441 O_4_4_1_3 WL_4_1 BL BLB W_4_4_3 W_4_4_3_bar CIM_cell
X3974 I441 O_4_4_1_4 WL_4_1 BL BLB W_4_4_4 W_4_4_4_bar CIM_cell
X3981 I442 O_4_4_2_1 WL_4_2 BL BLB W_4_4_1 W_4_4_1_bar CIM_cell
X3982 I442 O_4_4_2_2 WL_4_2 BL BLB W_4_4_2 W_4_4_2_bar CIM_cell
X3983 I442 O_4_4_2_3 WL_4_2 BL BLB W_4_4_3 W_4_4_3_bar CIM_cell
X3984 I442 O_4_4_2_4 WL_4_2 BL BLB W_4_4_4 W_4_4_4_bar CIM_cell
X3991 I443 O_4_4_3_1 WL_4_3 BL BLB W_4_4_1 W_4_4_1_bar CIM_cell
X3992 I443 O_4_4_3_2 WL_4_3 BL BLB W_4_4_2 W_4_4_2_bar CIM_cell
X3993 I443 O_4_4_3_3 WL_4_3 BL BLB W_4_4_3 W_4_4_3_bar CIM_cell
X3994 I443 O_4_4_3_4 WL_4_3 BL BLB W_4_4_4 W_4_4_4_bar CIM_cell
X4001 I444 O_4_4_4_1 WL_4_4 BL BLB W_4_4_1 W_4_4_1_bar CIM_cell
X4002 I444 O_4_4_4_2 WL_4_4 BL BLB W_4_4_2 W_4_4_2_bar CIM_cell
X4003 I444 O_4_4_4_3 WL_4_4 BL BLB W_4_4_3 W_4_4_3_bar CIM_cell
X4004 I444 O_4_4_4_4 WL_4_4 BL BLB W_4_4_4 W_4_4_4_bar CIM_cell
X4011 I451 O_4_5_1_1 WL_4_1 BL BLB W_4_5_1 W_4_5_1_bar CIM_cell
X4012 I451 O_4_5_1_2 WL_4_1 BL BLB W_4_5_2 W_4_5_2_bar CIM_cell
X4013 I451 O_4_5_1_3 WL_4_1 BL BLB W_4_5_3 W_4_5_3_bar CIM_cell
X4014 I451 O_4_5_1_4 WL_4_1 BL BLB W_4_5_4 W_4_5_4_bar CIM_cell
X4021 I452 O_4_5_2_1 WL_4_2 BL BLB W_4_5_1 W_4_5_1_bar CIM_cell
X4022 I452 O_4_5_2_2 WL_4_2 BL BLB W_4_5_2 W_4_5_2_bar CIM_cell
X4023 I452 O_4_5_2_3 WL_4_2 BL BLB W_4_5_3 W_4_5_3_bar CIM_cell
X4024 I452 O_4_5_2_4 WL_4_2 BL BLB W_4_5_4 W_4_5_4_bar CIM_cell
X4031 I453 O_4_5_3_1 WL_4_3 BL BLB W_4_5_1 W_4_5_1_bar CIM_cell
X4032 I453 O_4_5_3_2 WL_4_3 BL BLB W_4_5_2 W_4_5_2_bar CIM_cell
X4033 I453 O_4_5_3_3 WL_4_3 BL BLB W_4_5_3 W_4_5_3_bar CIM_cell
X4034 I453 O_4_5_3_4 WL_4_3 BL BLB W_4_5_4 W_4_5_4_bar CIM_cell
X4041 I454 O_4_5_4_1 WL_4_4 BL BLB W_4_5_1 W_4_5_1_bar CIM_cell
X4042 I454 O_4_5_4_2 WL_4_4 BL BLB W_4_5_2 W_4_5_2_bar CIM_cell
X4043 I454 O_4_5_4_3 WL_4_4 BL BLB W_4_5_3 W_4_5_3_bar CIM_cell
X4044 I454 O_4_5_4_4 WL_4_4 BL BLB W_4_5_4 W_4_5_4_bar CIM_cell
X4051 I461 O_4_6_1_1 WL_4_1 BL BLB W_4_6_1 W_4_6_1_bar CIM_cell
X4052 I461 O_4_6_1_2 WL_4_1 BL BLB W_4_6_2 W_4_6_2_bar CIM_cell
X4053 I461 O_4_6_1_3 WL_4_1 BL BLB W_4_6_3 W_4_6_3_bar CIM_cell
X4054 I461 O_4_6_1_4 WL_4_1 BL BLB W_4_6_4 W_4_6_4_bar CIM_cell
X4061 I462 O_4_6_2_1 WL_4_2 BL BLB W_4_6_1 W_4_6_1_bar CIM_cell
X4062 I462 O_4_6_2_2 WL_4_2 BL BLB W_4_6_2 W_4_6_2_bar CIM_cell
X4063 I462 O_4_6_2_3 WL_4_2 BL BLB W_4_6_3 W_4_6_3_bar CIM_cell
X4064 I462 O_4_6_2_4 WL_4_2 BL BLB W_4_6_4 W_4_6_4_bar CIM_cell
X4071 I463 O_4_6_3_1 WL_4_3 BL BLB W_4_6_1 W_4_6_1_bar CIM_cell
X4072 I463 O_4_6_3_2 WL_4_3 BL BLB W_4_6_2 W_4_6_2_bar CIM_cell
X4073 I463 O_4_6_3_3 WL_4_3 BL BLB W_4_6_3 W_4_6_3_bar CIM_cell
X4074 I463 O_4_6_3_4 WL_4_3 BL BLB W_4_6_4 W_4_6_4_bar CIM_cell
X4081 I464 O_4_6_4_1 WL_4_4 BL BLB W_4_6_1 W_4_6_1_bar CIM_cell
X4082 I464 O_4_6_4_2 WL_4_4 BL BLB W_4_6_2 W_4_6_2_bar CIM_cell
X4083 I464 O_4_6_4_3 WL_4_4 BL BLB W_4_6_3 W_4_6_3_bar CIM_cell
X4084 I464 O_4_6_4_4 WL_4_4 BL BLB W_4_6_4 W_4_6_4_bar CIM_cell
X4091 I471 O_4_7_1_1 WL_4_1 BL BLB W_4_7_1 W_4_7_1_bar CIM_cell
X4092 I471 O_4_7_1_2 WL_4_1 BL BLB W_4_7_2 W_4_7_2_bar CIM_cell
X4093 I471 O_4_7_1_3 WL_4_1 BL BLB W_4_7_3 W_4_7_3_bar CIM_cell
X4094 I471 O_4_7_1_4 WL_4_1 BL BLB W_4_7_4 W_4_7_4_bar CIM_cell
X4101 I472 O_4_7_2_1 WL_4_2 BL BLB W_4_7_1 W_4_7_1_bar CIM_cell
X4102 I472 O_4_7_2_2 WL_4_2 BL BLB W_4_7_2 W_4_7_2_bar CIM_cell
X4103 I472 O_4_7_2_3 WL_4_2 BL BLB W_4_7_3 W_4_7_3_bar CIM_cell
X4104 I472 O_4_7_2_4 WL_4_2 BL BLB W_4_7_4 W_4_7_4_bar CIM_cell
X4111 I473 O_4_7_3_1 WL_4_3 BL BLB W_4_7_1 W_4_7_1_bar CIM_cell
X4112 I473 O_4_7_3_2 WL_4_3 BL BLB W_4_7_2 W_4_7_2_bar CIM_cell
X4113 I473 O_4_7_3_3 WL_4_3 BL BLB W_4_7_3 W_4_7_3_bar CIM_cell
X4114 I473 O_4_7_3_4 WL_4_3 BL BLB W_4_7_4 W_4_7_4_bar CIM_cell
X4121 I474 O_4_7_4_1 WL_4_4 BL BLB W_4_7_1 W_4_7_1_bar CIM_cell
X4122 I474 O_4_7_4_2 WL_4_4 BL BLB W_4_7_2 W_4_7_2_bar CIM_cell
X4123 I474 O_4_7_4_3 WL_4_4 BL BLB W_4_7_3 W_4_7_3_bar CIM_cell
X4124 I474 O_4_7_4_4 WL_4_4 BL BLB W_4_7_4 W_4_7_4_bar CIM_cell
X4131 I481 O_4_8_1_1 WL_4_1 BL BLB W_4_8_1 W_4_8_1_bar CIM_cell
X4132 I481 O_4_8_1_2 WL_4_1 BL BLB W_4_8_2 W_4_8_2_bar CIM_cell
X4133 I481 O_4_8_1_3 WL_4_1 BL BLB W_4_8_3 W_4_8_3_bar CIM_cell
X4134 I481 O_4_8_1_4 WL_4_1 BL BLB W_4_8_4 W_4_8_4_bar CIM_cell
X4141 I482 O_4_8_2_1 WL_4_2 BL BLB W_4_8_1 W_4_8_1_bar CIM_cell
X4142 I482 O_4_8_2_2 WL_4_2 BL BLB W_4_8_2 W_4_8_2_bar CIM_cell
X4143 I482 O_4_8_2_3 WL_4_2 BL BLB W_4_8_3 W_4_8_3_bar CIM_cell
X4144 I482 O_4_8_2_4 WL_4_2 BL BLB W_4_8_4 W_4_8_4_bar CIM_cell
X4151 I483 O_4_8_3_1 WL_4_3 BL BLB W_4_8_1 W_4_8_1_bar CIM_cell
X4152 I483 O_4_8_3_2 WL_4_3 BL BLB W_4_8_2 W_4_8_2_bar CIM_cell
X4153 I483 O_4_8_3_3 WL_4_3 BL BLB W_4_8_3 W_4_8_3_bar CIM_cell
X4154 I483 O_4_8_3_4 WL_4_3 BL BLB W_4_8_4 W_4_8_4_bar CIM_cell
X4161 I484 O_4_8_4_1 WL_4_4 BL BLB W_4_8_1 W_4_8_1_bar CIM_cell
X4162 I484 O_4_8_4_2 WL_4_4 BL BLB W_4_8_2 W_4_8_2_bar CIM_cell
X4163 I484 O_4_8_4_3 WL_4_4 BL BLB W_4_8_3 W_4_8_3_bar CIM_cell
X4164 I484 O_4_8_4_4 WL_4_4 BL BLB W_4_8_4 W_4_8_4_bar CIM_cell
X4171 I491 O_4_9_1_1 WL_4_1 BL BLB W_4_9_1 W_4_9_1_bar CIM_cell
X4172 I491 O_4_9_1_2 WL_4_1 BL BLB W_4_9_2 W_4_9_2_bar CIM_cell
X4173 I491 O_4_9_1_3 WL_4_1 BL BLB W_4_9_3 W_4_9_3_bar CIM_cell
X4174 I491 O_4_9_1_4 WL_4_1 BL BLB W_4_9_4 W_4_9_4_bar CIM_cell
X4181 I492 O_4_9_2_1 WL_4_2 BL BLB W_4_9_1 W_4_9_1_bar CIM_cell
X4182 I492 O_4_9_2_2 WL_4_2 BL BLB W_4_9_2 W_4_9_2_bar CIM_cell
X4183 I492 O_4_9_2_3 WL_4_2 BL BLB W_4_9_3 W_4_9_3_bar CIM_cell
X4184 I492 O_4_9_2_4 WL_4_2 BL BLB W_4_9_4 W_4_9_4_bar CIM_cell
X4191 I493 O_4_9_3_1 WL_4_3 BL BLB W_4_9_1 W_4_9_1_bar CIM_cell
X4192 I493 O_4_9_3_2 WL_4_3 BL BLB W_4_9_2 W_4_9_2_bar CIM_cell
X4193 I493 O_4_9_3_3 WL_4_3 BL BLB W_4_9_3 W_4_9_3_bar CIM_cell
X4194 I493 O_4_9_3_4 WL_4_3 BL BLB W_4_9_4 W_4_9_4_bar CIM_cell
X4201 I494 O_4_9_4_1 WL_4_4 BL BLB W_4_9_1 W_4_9_1_bar CIM_cell
X4202 I494 O_4_9_4_2 WL_4_4 BL BLB W_4_9_2 W_4_9_2_bar CIM_cell
X4203 I494 O_4_9_4_3 WL_4_4 BL BLB W_4_9_3 W_4_9_3_bar CIM_cell
X4204 I494 O_4_9_4_4 WL_4_4 BL BLB W_4_9_4 W_4_9_4_bar CIM_cell
X4211 I4101 O_4_10_1_1 WL_4_1 BL BLB W_4_10_1 W_4_10_1_bar CIM_cell
X4212 I4101 O_4_10_1_2 WL_4_1 BL BLB W_4_10_2 W_4_10_2_bar CIM_cell
X4213 I4101 O_4_10_1_3 WL_4_1 BL BLB W_4_10_3 W_4_10_3_bar CIM_cell
X4214 I4101 O_4_10_1_4 WL_4_1 BL BLB W_4_10_4 W_4_10_4_bar CIM_cell
X4221 I4102 O_4_10_2_1 WL_4_2 BL BLB W_4_10_1 W_4_10_1_bar CIM_cell
X4222 I4102 O_4_10_2_2 WL_4_2 BL BLB W_4_10_2 W_4_10_2_bar CIM_cell
X4223 I4102 O_4_10_2_3 WL_4_2 BL BLB W_4_10_3 W_4_10_3_bar CIM_cell
X4224 I4102 O_4_10_2_4 WL_4_2 BL BLB W_4_10_4 W_4_10_4_bar CIM_cell
X4231 I4103 O_4_10_3_1 WL_4_3 BL BLB W_4_10_1 W_4_10_1_bar CIM_cell
X4232 I4103 O_4_10_3_2 WL_4_3 BL BLB W_4_10_2 W_4_10_2_bar CIM_cell
X4233 I4103 O_4_10_3_3 WL_4_3 BL BLB W_4_10_3 W_4_10_3_bar CIM_cell
X4234 I4103 O_4_10_3_4 WL_4_3 BL BLB W_4_10_4 W_4_10_4_bar CIM_cell
X4241 I4104 O_4_10_4_1 WL_4_4 BL BLB W_4_10_1 W_4_10_1_bar CIM_cell
X4242 I4104 O_4_10_4_2 WL_4_4 BL BLB W_4_10_2 W_4_10_2_bar CIM_cell
X4243 I4104 O_4_10_4_3 WL_4_4 BL BLB W_4_10_3 W_4_10_3_bar CIM_cell
X4244 I4104 O_4_10_4_4 WL_4_4 BL BLB W_4_10_4 W_4_10_4_bar CIM_cell
X4251 I4111 O_4_11_1_1 WL_4_1 BL BLB W_4_11_1 W_4_11_1_bar CIM_cell
X4252 I4111 O_4_11_1_2 WL_4_1 BL BLB W_4_11_2 W_4_11_2_bar CIM_cell
X4253 I4111 O_4_11_1_3 WL_4_1 BL BLB W_4_11_3 W_4_11_3_bar CIM_cell
X4254 I4111 O_4_11_1_4 WL_4_1 BL BLB W_4_11_4 W_4_11_4_bar CIM_cell
X4261 I4112 O_4_11_2_1 WL_4_2 BL BLB W_4_11_1 W_4_11_1_bar CIM_cell
X4262 I4112 O_4_11_2_2 WL_4_2 BL BLB W_4_11_2 W_4_11_2_bar CIM_cell
X4263 I4112 O_4_11_2_3 WL_4_2 BL BLB W_4_11_3 W_4_11_3_bar CIM_cell
X4264 I4112 O_4_11_2_4 WL_4_2 BL BLB W_4_11_4 W_4_11_4_bar CIM_cell
X4271 I4113 O_4_11_3_1 WL_4_3 BL BLB W_4_11_1 W_4_11_1_bar CIM_cell
X4272 I4113 O_4_11_3_2 WL_4_3 BL BLB W_4_11_2 W_4_11_2_bar CIM_cell
X4273 I4113 O_4_11_3_3 WL_4_3 BL BLB W_4_11_3 W_4_11_3_bar CIM_cell
X4274 I4113 O_4_11_3_4 WL_4_3 BL BLB W_4_11_4 W_4_11_4_bar CIM_cell
X4281 I4114 O_4_11_4_1 WL_4_4 BL BLB W_4_11_1 W_4_11_1_bar CIM_cell
X4282 I4114 O_4_11_4_2 WL_4_4 BL BLB W_4_11_2 W_4_11_2_bar CIM_cell
X4283 I4114 O_4_11_4_3 WL_4_4 BL BLB W_4_11_3 W_4_11_3_bar CIM_cell
X4284 I4114 O_4_11_4_4 WL_4_4 BL BLB W_4_11_4 W_4_11_4_bar CIM_cell
X4291 I4121 O_4_12_1_1 WL_4_1 BL BLB W_4_12_1 W_4_12_1_bar CIM_cell
X4292 I4121 O_4_12_1_2 WL_4_1 BL BLB W_4_12_2 W_4_12_2_bar CIM_cell
X4293 I4121 O_4_12_1_3 WL_4_1 BL BLB W_4_12_3 W_4_12_3_bar CIM_cell
X4294 I4121 O_4_12_1_4 WL_4_1 BL BLB W_4_12_4 W_4_12_4_bar CIM_cell
X4301 I4122 O_4_12_2_1 WL_4_2 BL BLB W_4_12_1 W_4_12_1_bar CIM_cell
X4302 I4122 O_4_12_2_2 WL_4_2 BL BLB W_4_12_2 W_4_12_2_bar CIM_cell
X4303 I4122 O_4_12_2_3 WL_4_2 BL BLB W_4_12_3 W_4_12_3_bar CIM_cell
X4304 I4122 O_4_12_2_4 WL_4_2 BL BLB W_4_12_4 W_4_12_4_bar CIM_cell
X4311 I4123 O_4_12_3_1 WL_4_3 BL BLB W_4_12_1 W_4_12_1_bar CIM_cell
X4312 I4123 O_4_12_3_2 WL_4_3 BL BLB W_4_12_2 W_4_12_2_bar CIM_cell
X4313 I4123 O_4_12_3_3 WL_4_3 BL BLB W_4_12_3 W_4_12_3_bar CIM_cell
X4314 I4123 O_4_12_3_4 WL_4_3 BL BLB W_4_12_4 W_4_12_4_bar CIM_cell
X4321 I4124 O_4_12_4_1 WL_4_4 BL BLB W_4_12_1 W_4_12_1_bar CIM_cell
X4322 I4124 O_4_12_4_2 WL_4_4 BL BLB W_4_12_2 W_4_12_2_bar CIM_cell
X4323 I4124 O_4_12_4_3 WL_4_4 BL BLB W_4_12_3 W_4_12_3_bar CIM_cell
X4324 I4124 O_4_12_4_4 WL_4_4 BL BLB W_4_12_4 W_4_12_4_bar CIM_cell
X4331 I4131 O_4_13_1_1 WL_4_1 BL BLB W_4_13_1 W_4_13_1_bar CIM_cell
X4332 I4131 O_4_13_1_2 WL_4_1 BL BLB W_4_13_2 W_4_13_2_bar CIM_cell
X4333 I4131 O_4_13_1_3 WL_4_1 BL BLB W_4_13_3 W_4_13_3_bar CIM_cell
X4334 I4131 O_4_13_1_4 WL_4_1 BL BLB W_4_13_4 W_4_13_4_bar CIM_cell
X4341 I4132 O_4_13_2_1 WL_4_2 BL BLB W_4_13_1 W_4_13_1_bar CIM_cell
X4342 I4132 O_4_13_2_2 WL_4_2 BL BLB W_4_13_2 W_4_13_2_bar CIM_cell
X4343 I4132 O_4_13_2_3 WL_4_2 BL BLB W_4_13_3 W_4_13_3_bar CIM_cell
X4344 I4132 O_4_13_2_4 WL_4_2 BL BLB W_4_13_4 W_4_13_4_bar CIM_cell
X4351 I4133 O_4_13_3_1 WL_4_3 BL BLB W_4_13_1 W_4_13_1_bar CIM_cell
X4352 I4133 O_4_13_3_2 WL_4_3 BL BLB W_4_13_2 W_4_13_2_bar CIM_cell
X4353 I4133 O_4_13_3_3 WL_4_3 BL BLB W_4_13_3 W_4_13_3_bar CIM_cell
X4354 I4133 O_4_13_3_4 WL_4_3 BL BLB W_4_13_4 W_4_13_4_bar CIM_cell
X4361 I4134 O_4_13_4_1 WL_4_4 BL BLB W_4_13_1 W_4_13_1_bar CIM_cell
X4362 I4134 O_4_13_4_2 WL_4_4 BL BLB W_4_13_2 W_4_13_2_bar CIM_cell
X4363 I4134 O_4_13_4_3 WL_4_4 BL BLB W_4_13_3 W_4_13_3_bar CIM_cell
X4364 I4134 O_4_13_4_4 WL_4_4 BL BLB W_4_13_4 W_4_13_4_bar CIM_cell
X4371 I4141 O_4_14_1_1 WL_4_1 BL BLB W_4_14_1 W_4_14_1_bar CIM_cell
X4372 I4141 O_4_14_1_2 WL_4_1 BL BLB W_4_14_2 W_4_14_2_bar CIM_cell
X4373 I4141 O_4_14_1_3 WL_4_1 BL BLB W_4_14_3 W_4_14_3_bar CIM_cell
X4374 I4141 O_4_14_1_4 WL_4_1 BL BLB W_4_14_4 W_4_14_4_bar CIM_cell
X4381 I4142 O_4_14_2_1 WL_4_2 BL BLB W_4_14_1 W_4_14_1_bar CIM_cell
X4382 I4142 O_4_14_2_2 WL_4_2 BL BLB W_4_14_2 W_4_14_2_bar CIM_cell
X4383 I4142 O_4_14_2_3 WL_4_2 BL BLB W_4_14_3 W_4_14_3_bar CIM_cell
X4384 I4142 O_4_14_2_4 WL_4_2 BL BLB W_4_14_4 W_4_14_4_bar CIM_cell
X4391 I4143 O_4_14_3_1 WL_4_3 BL BLB W_4_14_1 W_4_14_1_bar CIM_cell
X4392 I4143 O_4_14_3_2 WL_4_3 BL BLB W_4_14_2 W_4_14_2_bar CIM_cell
X4393 I4143 O_4_14_3_3 WL_4_3 BL BLB W_4_14_3 W_4_14_3_bar CIM_cell
X4394 I4143 O_4_14_3_4 WL_4_3 BL BLB W_4_14_4 W_4_14_4_bar CIM_cell
X4401 I4144 O_4_14_4_1 WL_4_4 BL BLB W_4_14_1 W_4_14_1_bar CIM_cell
X4402 I4144 O_4_14_4_2 WL_4_4 BL BLB W_4_14_2 W_4_14_2_bar CIM_cell
X4403 I4144 O_4_14_4_3 WL_4_4 BL BLB W_4_14_3 W_4_14_3_bar CIM_cell
X4404 I4144 O_4_14_4_4 WL_4_4 BL BLB W_4_14_4 W_4_14_4_bar CIM_cell
X4411 I4151 O_4_15_1_1 WL_4_1 BL BLB W_4_15_1 W_4_15_1_bar CIM_cell
X4412 I4151 O_4_15_1_2 WL_4_1 BL BLB W_4_15_2 W_4_15_2_bar CIM_cell
X4413 I4151 O_4_15_1_3 WL_4_1 BL BLB W_4_15_3 W_4_15_3_bar CIM_cell
X4414 I4151 O_4_15_1_4 WL_4_1 BL BLB W_4_15_4 W_4_15_4_bar CIM_cell
X4421 I4152 O_4_15_2_1 WL_4_2 BL BLB W_4_15_1 W_4_15_1_bar CIM_cell
X4422 I4152 O_4_15_2_2 WL_4_2 BL BLB W_4_15_2 W_4_15_2_bar CIM_cell
X4423 I4152 O_4_15_2_3 WL_4_2 BL BLB W_4_15_3 W_4_15_3_bar CIM_cell
X4424 I4152 O_4_15_2_4 WL_4_2 BL BLB W_4_15_4 W_4_15_4_bar CIM_cell
X4431 I4153 O_4_15_3_1 WL_4_3 BL BLB W_4_15_1 W_4_15_1_bar CIM_cell
X4432 I4153 O_4_15_3_2 WL_4_3 BL BLB W_4_15_2 W_4_15_2_bar CIM_cell
X4433 I4153 O_4_15_3_3 WL_4_3 BL BLB W_4_15_3 W_4_15_3_bar CIM_cell
X4434 I4153 O_4_15_3_4 WL_4_3 BL BLB W_4_15_4 W_4_15_4_bar CIM_cell
X4441 I4154 O_4_15_4_1 WL_4_4 BL BLB W_4_15_1 W_4_15_1_bar CIM_cell
X4442 I4154 O_4_15_4_2 WL_4_4 BL BLB W_4_15_2 W_4_15_2_bar CIM_cell
X4443 I4154 O_4_15_4_3 WL_4_4 BL BLB W_4_15_3 W_4_15_3_bar CIM_cell
X4444 I4154 O_4_15_4_4 WL_4_4 BL BLB W_4_15_4 W_4_15_4_bar CIM_cell
X4451 I4161 O_4_16_1_1 WL_4_1 BL BLB W_4_16_1 W_4_16_1_bar CIM_cell
X4452 I4161 O_4_16_1_2 WL_4_1 BL BLB W_4_16_2 W_4_16_2_bar CIM_cell
X4453 I4161 O_4_16_1_3 WL_4_1 BL BLB W_4_16_3 W_4_16_3_bar CIM_cell
X4454 I4161 O_4_16_1_4 WL_4_1 BL BLB W_4_16_4 W_4_16_4_bar CIM_cell
X4461 I4162 O_4_16_2_1 WL_4_2 BL BLB W_4_16_1 W_4_16_1_bar CIM_cell
X4462 I4162 O_4_16_2_2 WL_4_2 BL BLB W_4_16_2 W_4_16_2_bar CIM_cell
X4463 I4162 O_4_16_2_3 WL_4_2 BL BLB W_4_16_3 W_4_16_3_bar CIM_cell
X4464 I4162 O_4_16_2_4 WL_4_2 BL BLB W_4_16_4 W_4_16_4_bar CIM_cell
X4471 I4163 O_4_16_3_1 WL_4_3 BL BLB W_4_16_1 W_4_16_1_bar CIM_cell
X4472 I4163 O_4_16_3_2 WL_4_3 BL BLB W_4_16_2 W_4_16_2_bar CIM_cell
X4473 I4163 O_4_16_3_3 WL_4_3 BL BLB W_4_16_3 W_4_16_3_bar CIM_cell
X4474 I4163 O_4_16_3_4 WL_4_3 BL BLB W_4_16_4 W_4_16_4_bar CIM_cell
X4481 I4164 O_4_16_4_1 WL_4_4 BL BLB W_4_16_1 W_4_16_1_bar CIM_cell
X4482 I4164 O_4_16_4_2 WL_4_4 BL BLB W_4_16_2 W_4_16_2_bar CIM_cell
X4483 I4164 O_4_16_4_3 WL_4_4 BL BLB W_4_16_3 W_4_16_3_bar CIM_cell
X4484 I4164 O_4_16_4_4 WL_4_4 BL BLB W_4_16_4 W_4_16_4_bar CIM_cell
X4491 I4171 O_4_17_1_1 WL_4_1 BL BLB W_4_17_1 W_4_17_1_bar CIM_cell
X4492 I4171 O_4_17_1_2 WL_4_1 BL BLB W_4_17_2 W_4_17_2_bar CIM_cell
X4493 I4171 O_4_17_1_3 WL_4_1 BL BLB W_4_17_3 W_4_17_3_bar CIM_cell
X4494 I4171 O_4_17_1_4 WL_4_1 BL BLB W_4_17_4 W_4_17_4_bar CIM_cell
X4501 I4172 O_4_17_2_1 WL_4_2 BL BLB W_4_17_1 W_4_17_1_bar CIM_cell
X4502 I4172 O_4_17_2_2 WL_4_2 BL BLB W_4_17_2 W_4_17_2_bar CIM_cell
X4503 I4172 O_4_17_2_3 WL_4_2 BL BLB W_4_17_3 W_4_17_3_bar CIM_cell
X4504 I4172 O_4_17_2_4 WL_4_2 BL BLB W_4_17_4 W_4_17_4_bar CIM_cell
X4511 I4173 O_4_17_3_1 WL_4_3 BL BLB W_4_17_1 W_4_17_1_bar CIM_cell
X4512 I4173 O_4_17_3_2 WL_4_3 BL BLB W_4_17_2 W_4_17_2_bar CIM_cell
X4513 I4173 O_4_17_3_3 WL_4_3 BL BLB W_4_17_3 W_4_17_3_bar CIM_cell
X4514 I4173 O_4_17_3_4 WL_4_3 BL BLB W_4_17_4 W_4_17_4_bar CIM_cell
X4521 I4174 O_4_17_4_1 WL_4_4 BL BLB W_4_17_1 W_4_17_1_bar CIM_cell
X4522 I4174 O_4_17_4_2 WL_4_4 BL BLB W_4_17_2 W_4_17_2_bar CIM_cell
X4523 I4174 O_4_17_4_3 WL_4_4 BL BLB W_4_17_3 W_4_17_3_bar CIM_cell
X4524 I4174 O_4_17_4_4 WL_4_4 BL BLB W_4_17_4 W_4_17_4_bar CIM_cell
X4531 I4181 O_4_18_1_1 WL_4_1 BL BLB W_4_18_1 W_4_18_1_bar CIM_cell
X4532 I4181 O_4_18_1_2 WL_4_1 BL BLB W_4_18_2 W_4_18_2_bar CIM_cell
X4533 I4181 O_4_18_1_3 WL_4_1 BL BLB W_4_18_3 W_4_18_3_bar CIM_cell
X4534 I4181 O_4_18_1_4 WL_4_1 BL BLB W_4_18_4 W_4_18_4_bar CIM_cell
X4541 I4182 O_4_18_2_1 WL_4_2 BL BLB W_4_18_1 W_4_18_1_bar CIM_cell
X4542 I4182 O_4_18_2_2 WL_4_2 BL BLB W_4_18_2 W_4_18_2_bar CIM_cell
X4543 I4182 O_4_18_2_3 WL_4_2 BL BLB W_4_18_3 W_4_18_3_bar CIM_cell
X4544 I4182 O_4_18_2_4 WL_4_2 BL BLB W_4_18_4 W_4_18_4_bar CIM_cell
X4551 I4183 O_4_18_3_1 WL_4_3 BL BLB W_4_18_1 W_4_18_1_bar CIM_cell
X4552 I4183 O_4_18_3_2 WL_4_3 BL BLB W_4_18_2 W_4_18_2_bar CIM_cell
X4553 I4183 O_4_18_3_3 WL_4_3 BL BLB W_4_18_3 W_4_18_3_bar CIM_cell
X4554 I4183 O_4_18_3_4 WL_4_3 BL BLB W_4_18_4 W_4_18_4_bar CIM_cell
X4561 I4184 O_4_18_4_1 WL_4_4 BL BLB W_4_18_1 W_4_18_1_bar CIM_cell
X4562 I4184 O_4_18_4_2 WL_4_4 BL BLB W_4_18_2 W_4_18_2_bar CIM_cell
X4563 I4184 O_4_18_4_3 WL_4_4 BL BLB W_4_18_3 W_4_18_3_bar CIM_cell
X4564 I4184 O_4_18_4_4 WL_4_4 BL BLB W_4_18_4 W_4_18_4_bar CIM_cell
X4571 I4191 O_4_19_1_1 WL_4_1 BL BLB W_4_19_1 W_4_19_1_bar CIM_cell
X4572 I4191 O_4_19_1_2 WL_4_1 BL BLB W_4_19_2 W_4_19_2_bar CIM_cell
X4573 I4191 O_4_19_1_3 WL_4_1 BL BLB W_4_19_3 W_4_19_3_bar CIM_cell
X4574 I4191 O_4_19_1_4 WL_4_1 BL BLB W_4_19_4 W_4_19_4_bar CIM_cell
X4581 I4192 O_4_19_2_1 WL_4_2 BL BLB W_4_19_1 W_4_19_1_bar CIM_cell
X4582 I4192 O_4_19_2_2 WL_4_2 BL BLB W_4_19_2 W_4_19_2_bar CIM_cell
X4583 I4192 O_4_19_2_3 WL_4_2 BL BLB W_4_19_3 W_4_19_3_bar CIM_cell
X4584 I4192 O_4_19_2_4 WL_4_2 BL BLB W_4_19_4 W_4_19_4_bar CIM_cell
X4591 I4193 O_4_19_3_1 WL_4_3 BL BLB W_4_19_1 W_4_19_1_bar CIM_cell
X4592 I4193 O_4_19_3_2 WL_4_3 BL BLB W_4_19_2 W_4_19_2_bar CIM_cell
X4593 I4193 O_4_19_3_3 WL_4_3 BL BLB W_4_19_3 W_4_19_3_bar CIM_cell
X4594 I4193 O_4_19_3_4 WL_4_3 BL BLB W_4_19_4 W_4_19_4_bar CIM_cell
X4601 I4194 O_4_19_4_1 WL_4_4 BL BLB W_4_19_1 W_4_19_1_bar CIM_cell
X4602 I4194 O_4_19_4_2 WL_4_4 BL BLB W_4_19_2 W_4_19_2_bar CIM_cell
X4603 I4194 O_4_19_4_3 WL_4_4 BL BLB W_4_19_3 W_4_19_3_bar CIM_cell
X4604 I4194 O_4_19_4_4 WL_4_4 BL BLB W_4_19_4 W_4_19_4_bar CIM_cell
X4611 I4201 O_4_20_1_1 WL_4_1 BL BLB W_4_20_1 W_4_20_1_bar CIM_cell
X4612 I4201 O_4_20_1_2 WL_4_1 BL BLB W_4_20_2 W_4_20_2_bar CIM_cell
X4613 I4201 O_4_20_1_3 WL_4_1 BL BLB W_4_20_3 W_4_20_3_bar CIM_cell
X4614 I4201 O_4_20_1_4 WL_4_1 BL BLB W_4_20_4 W_4_20_4_bar CIM_cell
X4621 I4202 O_4_20_2_1 WL_4_2 BL BLB W_4_20_1 W_4_20_1_bar CIM_cell
X4622 I4202 O_4_20_2_2 WL_4_2 BL BLB W_4_20_2 W_4_20_2_bar CIM_cell
X4623 I4202 O_4_20_2_3 WL_4_2 BL BLB W_4_20_3 W_4_20_3_bar CIM_cell
X4624 I4202 O_4_20_2_4 WL_4_2 BL BLB W_4_20_4 W_4_20_4_bar CIM_cell
X4631 I4203 O_4_20_3_1 WL_4_3 BL BLB W_4_20_1 W_4_20_1_bar CIM_cell
X4632 I4203 O_4_20_3_2 WL_4_3 BL BLB W_4_20_2 W_4_20_2_bar CIM_cell
X4633 I4203 O_4_20_3_3 WL_4_3 BL BLB W_4_20_3 W_4_20_3_bar CIM_cell
X4634 I4203 O_4_20_3_4 WL_4_3 BL BLB W_4_20_4 W_4_20_4_bar CIM_cell
X4641 I4204 O_4_20_4_1 WL_4_4 BL BLB W_4_20_1 W_4_20_1_bar CIM_cell
X4642 I4204 O_4_20_4_2 WL_4_4 BL BLB W_4_20_2 W_4_20_2_bar CIM_cell
X4643 I4204 O_4_20_4_3 WL_4_4 BL BLB W_4_20_3 W_4_20_3_bar CIM_cell
X4644 I4204 O_4_20_4_4 WL_4_4 BL BLB W_4_20_4 W_4_20_4_bar CIM_cell
X4651 I4211 O_4_21_1_1 WL_4_1 BL BLB W_4_21_1 W_4_21_1_bar CIM_cell
X4652 I4211 O_4_21_1_2 WL_4_1 BL BLB W_4_21_2 W_4_21_2_bar CIM_cell
X4653 I4211 O_4_21_1_3 WL_4_1 BL BLB W_4_21_3 W_4_21_3_bar CIM_cell
X4654 I4211 O_4_21_1_4 WL_4_1 BL BLB W_4_21_4 W_4_21_4_bar CIM_cell
X4661 I4212 O_4_21_2_1 WL_4_2 BL BLB W_4_21_1 W_4_21_1_bar CIM_cell
X4662 I4212 O_4_21_2_2 WL_4_2 BL BLB W_4_21_2 W_4_21_2_bar CIM_cell
X4663 I4212 O_4_21_2_3 WL_4_2 BL BLB W_4_21_3 W_4_21_3_bar CIM_cell
X4664 I4212 O_4_21_2_4 WL_4_2 BL BLB W_4_21_4 W_4_21_4_bar CIM_cell
X4671 I4213 O_4_21_3_1 WL_4_3 BL BLB W_4_21_1 W_4_21_1_bar CIM_cell
X4672 I4213 O_4_21_3_2 WL_4_3 BL BLB W_4_21_2 W_4_21_2_bar CIM_cell
X4673 I4213 O_4_21_3_3 WL_4_3 BL BLB W_4_21_3 W_4_21_3_bar CIM_cell
X4674 I4213 O_4_21_3_4 WL_4_3 BL BLB W_4_21_4 W_4_21_4_bar CIM_cell
X4681 I4214 O_4_21_4_1 WL_4_4 BL BLB W_4_21_1 W_4_21_1_bar CIM_cell
X4682 I4214 O_4_21_4_2 WL_4_4 BL BLB W_4_21_2 W_4_21_2_bar CIM_cell
X4683 I4214 O_4_21_4_3 WL_4_4 BL BLB W_4_21_3 W_4_21_3_bar CIM_cell
X4684 I4214 O_4_21_4_4 WL_4_4 BL BLB W_4_21_4 W_4_21_4_bar CIM_cell
X4691 I4221 O_4_22_1_1 WL_4_1 BL BLB W_4_22_1 W_4_22_1_bar CIM_cell
X4692 I4221 O_4_22_1_2 WL_4_1 BL BLB W_4_22_2 W_4_22_2_bar CIM_cell
X4693 I4221 O_4_22_1_3 WL_4_1 BL BLB W_4_22_3 W_4_22_3_bar CIM_cell
X4694 I4221 O_4_22_1_4 WL_4_1 BL BLB W_4_22_4 W_4_22_4_bar CIM_cell
X4701 I4222 O_4_22_2_1 WL_4_2 BL BLB W_4_22_1 W_4_22_1_bar CIM_cell
X4702 I4222 O_4_22_2_2 WL_4_2 BL BLB W_4_22_2 W_4_22_2_bar CIM_cell
X4703 I4222 O_4_22_2_3 WL_4_2 BL BLB W_4_22_3 W_4_22_3_bar CIM_cell
X4704 I4222 O_4_22_2_4 WL_4_2 BL BLB W_4_22_4 W_4_22_4_bar CIM_cell
X4711 I4223 O_4_22_3_1 WL_4_3 BL BLB W_4_22_1 W_4_22_1_bar CIM_cell
X4712 I4223 O_4_22_3_2 WL_4_3 BL BLB W_4_22_2 W_4_22_2_bar CIM_cell
X4713 I4223 O_4_22_3_3 WL_4_3 BL BLB W_4_22_3 W_4_22_3_bar CIM_cell
X4714 I4223 O_4_22_3_4 WL_4_3 BL BLB W_4_22_4 W_4_22_4_bar CIM_cell
X4721 I4224 O_4_22_4_1 WL_4_4 BL BLB W_4_22_1 W_4_22_1_bar CIM_cell
X4722 I4224 O_4_22_4_2 WL_4_4 BL BLB W_4_22_2 W_4_22_2_bar CIM_cell
X4723 I4224 O_4_22_4_3 WL_4_4 BL BLB W_4_22_3 W_4_22_3_bar CIM_cell
X4724 I4224 O_4_22_4_4 WL_4_4 BL BLB W_4_22_4 W_4_22_4_bar CIM_cell
X4731 I4231 O_4_23_1_1 WL_4_1 BL BLB W_4_23_1 W_4_23_1_bar CIM_cell
X4732 I4231 O_4_23_1_2 WL_4_1 BL BLB W_4_23_2 W_4_23_2_bar CIM_cell
X4733 I4231 O_4_23_1_3 WL_4_1 BL BLB W_4_23_3 W_4_23_3_bar CIM_cell
X4734 I4231 O_4_23_1_4 WL_4_1 BL BLB W_4_23_4 W_4_23_4_bar CIM_cell
X4741 I4232 O_4_23_2_1 WL_4_2 BL BLB W_4_23_1 W_4_23_1_bar CIM_cell
X4742 I4232 O_4_23_2_2 WL_4_2 BL BLB W_4_23_2 W_4_23_2_bar CIM_cell
X4743 I4232 O_4_23_2_3 WL_4_2 BL BLB W_4_23_3 W_4_23_3_bar CIM_cell
X4744 I4232 O_4_23_2_4 WL_4_2 BL BLB W_4_23_4 W_4_23_4_bar CIM_cell
X4751 I4233 O_4_23_3_1 WL_4_3 BL BLB W_4_23_1 W_4_23_1_bar CIM_cell
X4752 I4233 O_4_23_3_2 WL_4_3 BL BLB W_4_23_2 W_4_23_2_bar CIM_cell
X4753 I4233 O_4_23_3_3 WL_4_3 BL BLB W_4_23_3 W_4_23_3_bar CIM_cell
X4754 I4233 O_4_23_3_4 WL_4_3 BL BLB W_4_23_4 W_4_23_4_bar CIM_cell
X4761 I4234 O_4_23_4_1 WL_4_4 BL BLB W_4_23_1 W_4_23_1_bar CIM_cell
X4762 I4234 O_4_23_4_2 WL_4_4 BL BLB W_4_23_2 W_4_23_2_bar CIM_cell
X4763 I4234 O_4_23_4_3 WL_4_4 BL BLB W_4_23_3 W_4_23_3_bar CIM_cell
X4764 I4234 O_4_23_4_4 WL_4_4 BL BLB W_4_23_4 W_4_23_4_bar CIM_cell
X4771 I4241 O_4_24_1_1 WL_4_1 BL BLB W_4_24_1 W_4_24_1_bar CIM_cell
X4772 I4241 O_4_24_1_2 WL_4_1 BL BLB W_4_24_2 W_4_24_2_bar CIM_cell
X4773 I4241 O_4_24_1_3 WL_4_1 BL BLB W_4_24_3 W_4_24_3_bar CIM_cell
X4774 I4241 O_4_24_1_4 WL_4_1 BL BLB W_4_24_4 W_4_24_4_bar CIM_cell
X4781 I4242 O_4_24_2_1 WL_4_2 BL BLB W_4_24_1 W_4_24_1_bar CIM_cell
X4782 I4242 O_4_24_2_2 WL_4_2 BL BLB W_4_24_2 W_4_24_2_bar CIM_cell
X4783 I4242 O_4_24_2_3 WL_4_2 BL BLB W_4_24_3 W_4_24_3_bar CIM_cell
X4784 I4242 O_4_24_2_4 WL_4_2 BL BLB W_4_24_4 W_4_24_4_bar CIM_cell
X4791 I4243 O_4_24_3_1 WL_4_3 BL BLB W_4_24_1 W_4_24_1_bar CIM_cell
X4792 I4243 O_4_24_3_2 WL_4_3 BL BLB W_4_24_2 W_4_24_2_bar CIM_cell
X4793 I4243 O_4_24_3_3 WL_4_3 BL BLB W_4_24_3 W_4_24_3_bar CIM_cell
X4794 I4243 O_4_24_3_4 WL_4_3 BL BLB W_4_24_4 W_4_24_4_bar CIM_cell
X4801 I4244 O_4_24_4_1 WL_4_4 BL BLB W_4_24_1 W_4_24_1_bar CIM_cell
X4802 I4244 O_4_24_4_2 WL_4_4 BL BLB W_4_24_2 W_4_24_2_bar CIM_cell
X4803 I4244 O_4_24_4_3 WL_4_4 BL BLB W_4_24_3 W_4_24_3_bar CIM_cell
X4804 I4244 O_4_24_4_4 WL_4_4 BL BLB W_4_24_4 W_4_24_4_bar CIM_cell
X4811 I4251 O_4_25_1_1 WL_4_1 BL BLB W_4_25_1 W_4_25_1_bar CIM_cell
X4812 I4251 O_4_25_1_2 WL_4_1 BL BLB W_4_25_2 W_4_25_2_bar CIM_cell
X4813 I4251 O_4_25_1_3 WL_4_1 BL BLB W_4_25_3 W_4_25_3_bar CIM_cell
X4814 I4251 O_4_25_1_4 WL_4_1 BL BLB W_4_25_4 W_4_25_4_bar CIM_cell
X4821 I4252 O_4_25_2_1 WL_4_2 BL BLB W_4_25_1 W_4_25_1_bar CIM_cell
X4822 I4252 O_4_25_2_2 WL_4_2 BL BLB W_4_25_2 W_4_25_2_bar CIM_cell
X4823 I4252 O_4_25_2_3 WL_4_2 BL BLB W_4_25_3 W_4_25_3_bar CIM_cell
X4824 I4252 O_4_25_2_4 WL_4_2 BL BLB W_4_25_4 W_4_25_4_bar CIM_cell
X4831 I4253 O_4_25_3_1 WL_4_3 BL BLB W_4_25_1 W_4_25_1_bar CIM_cell
X4832 I4253 O_4_25_3_2 WL_4_3 BL BLB W_4_25_2 W_4_25_2_bar CIM_cell
X4833 I4253 O_4_25_3_3 WL_4_3 BL BLB W_4_25_3 W_4_25_3_bar CIM_cell
X4834 I4253 O_4_25_3_4 WL_4_3 BL BLB W_4_25_4 W_4_25_4_bar CIM_cell
X4841 I4254 O_4_25_4_1 WL_4_4 BL BLB W_4_25_1 W_4_25_1_bar CIM_cell
X4842 I4254 O_4_25_4_2 WL_4_4 BL BLB W_4_25_2 W_4_25_2_bar CIM_cell
X4843 I4254 O_4_25_4_3 WL_4_4 BL BLB W_4_25_3 W_4_25_3_bar CIM_cell
X4844 I4254 O_4_25_4_4 WL_4_4 BL BLB W_4_25_4 W_4_25_4_bar CIM_cell
X4851 I4261 O_4_26_1_1 WL_4_1 BL BLB W_4_26_1 W_4_26_1_bar CIM_cell
X4852 I4261 O_4_26_1_2 WL_4_1 BL BLB W_4_26_2 W_4_26_2_bar CIM_cell
X4853 I4261 O_4_26_1_3 WL_4_1 BL BLB W_4_26_3 W_4_26_3_bar CIM_cell
X4854 I4261 O_4_26_1_4 WL_4_1 BL BLB W_4_26_4 W_4_26_4_bar CIM_cell
X4861 I4262 O_4_26_2_1 WL_4_2 BL BLB W_4_26_1 W_4_26_1_bar CIM_cell
X4862 I4262 O_4_26_2_2 WL_4_2 BL BLB W_4_26_2 W_4_26_2_bar CIM_cell
X4863 I4262 O_4_26_2_3 WL_4_2 BL BLB W_4_26_3 W_4_26_3_bar CIM_cell
X4864 I4262 O_4_26_2_4 WL_4_2 BL BLB W_4_26_4 W_4_26_4_bar CIM_cell
X4871 I4263 O_4_26_3_1 WL_4_3 BL BLB W_4_26_1 W_4_26_1_bar CIM_cell
X4872 I4263 O_4_26_3_2 WL_4_3 BL BLB W_4_26_2 W_4_26_2_bar CIM_cell
X4873 I4263 O_4_26_3_3 WL_4_3 BL BLB W_4_26_3 W_4_26_3_bar CIM_cell
X4874 I4263 O_4_26_3_4 WL_4_3 BL BLB W_4_26_4 W_4_26_4_bar CIM_cell
X4881 I4264 O_4_26_4_1 WL_4_4 BL BLB W_4_26_1 W_4_26_1_bar CIM_cell
X4882 I4264 O_4_26_4_2 WL_4_4 BL BLB W_4_26_2 W_4_26_2_bar CIM_cell
X4883 I4264 O_4_26_4_3 WL_4_4 BL BLB W_4_26_3 W_4_26_3_bar CIM_cell
X4884 I4264 O_4_26_4_4 WL_4_4 BL BLB W_4_26_4 W_4_26_4_bar CIM_cell
X4891 I4271 O_4_27_1_1 WL_4_1 BL BLB W_4_27_1 W_4_27_1_bar CIM_cell
X4892 I4271 O_4_27_1_2 WL_4_1 BL BLB W_4_27_2 W_4_27_2_bar CIM_cell
X4893 I4271 O_4_27_1_3 WL_4_1 BL BLB W_4_27_3 W_4_27_3_bar CIM_cell
X4894 I4271 O_4_27_1_4 WL_4_1 BL BLB W_4_27_4 W_4_27_4_bar CIM_cell
X4901 I4272 O_4_27_2_1 WL_4_2 BL BLB W_4_27_1 W_4_27_1_bar CIM_cell
X4902 I4272 O_4_27_2_2 WL_4_2 BL BLB W_4_27_2 W_4_27_2_bar CIM_cell
X4903 I4272 O_4_27_2_3 WL_4_2 BL BLB W_4_27_3 W_4_27_3_bar CIM_cell
X4904 I4272 O_4_27_2_4 WL_4_2 BL BLB W_4_27_4 W_4_27_4_bar CIM_cell
X4911 I4273 O_4_27_3_1 WL_4_3 BL BLB W_4_27_1 W_4_27_1_bar CIM_cell
X4912 I4273 O_4_27_3_2 WL_4_3 BL BLB W_4_27_2 W_4_27_2_bar CIM_cell
X4913 I4273 O_4_27_3_3 WL_4_3 BL BLB W_4_27_3 W_4_27_3_bar CIM_cell
X4914 I4273 O_4_27_3_4 WL_4_3 BL BLB W_4_27_4 W_4_27_4_bar CIM_cell
X4921 I4274 O_4_27_4_1 WL_4_4 BL BLB W_4_27_1 W_4_27_1_bar CIM_cell
X4922 I4274 O_4_27_4_2 WL_4_4 BL BLB W_4_27_2 W_4_27_2_bar CIM_cell
X4923 I4274 O_4_27_4_3 WL_4_4 BL BLB W_4_27_3 W_4_27_3_bar CIM_cell
X4924 I4274 O_4_27_4_4 WL_4_4 BL BLB W_4_27_4 W_4_27_4_bar CIM_cell
X4931 I4281 O_4_28_1_1 WL_4_1 BL BLB W_4_28_1 W_4_28_1_bar CIM_cell
X4932 I4281 O_4_28_1_2 WL_4_1 BL BLB W_4_28_2 W_4_28_2_bar CIM_cell
X4933 I4281 O_4_28_1_3 WL_4_1 BL BLB W_4_28_3 W_4_28_3_bar CIM_cell
X4934 I4281 O_4_28_1_4 WL_4_1 BL BLB W_4_28_4 W_4_28_4_bar CIM_cell
X4941 I4282 O_4_28_2_1 WL_4_2 BL BLB W_4_28_1 W_4_28_1_bar CIM_cell
X4942 I4282 O_4_28_2_2 WL_4_2 BL BLB W_4_28_2 W_4_28_2_bar CIM_cell
X4943 I4282 O_4_28_2_3 WL_4_2 BL BLB W_4_28_3 W_4_28_3_bar CIM_cell
X4944 I4282 O_4_28_2_4 WL_4_2 BL BLB W_4_28_4 W_4_28_4_bar CIM_cell
X4951 I4283 O_4_28_3_1 WL_4_3 BL BLB W_4_28_1 W_4_28_1_bar CIM_cell
X4952 I4283 O_4_28_3_2 WL_4_3 BL BLB W_4_28_2 W_4_28_2_bar CIM_cell
X4953 I4283 O_4_28_3_3 WL_4_3 BL BLB W_4_28_3 W_4_28_3_bar CIM_cell
X4954 I4283 O_4_28_3_4 WL_4_3 BL BLB W_4_28_4 W_4_28_4_bar CIM_cell
X4961 I4284 O_4_28_4_1 WL_4_4 BL BLB W_4_28_1 W_4_28_1_bar CIM_cell
X4962 I4284 O_4_28_4_2 WL_4_4 BL BLB W_4_28_2 W_4_28_2_bar CIM_cell
X4963 I4284 O_4_28_4_3 WL_4_4 BL BLB W_4_28_3 W_4_28_3_bar CIM_cell
X4964 I4284 O_4_28_4_4 WL_4_4 BL BLB W_4_28_4 W_4_28_4_bar CIM_cell
X4971 I4291 O_4_29_1_1 WL_4_1 BL BLB W_4_29_1 W_4_29_1_bar CIM_cell
X4972 I4291 O_4_29_1_2 WL_4_1 BL BLB W_4_29_2 W_4_29_2_bar CIM_cell
X4973 I4291 O_4_29_1_3 WL_4_1 BL BLB W_4_29_3 W_4_29_3_bar CIM_cell
X4974 I4291 O_4_29_1_4 WL_4_1 BL BLB W_4_29_4 W_4_29_4_bar CIM_cell
X4981 I4292 O_4_29_2_1 WL_4_2 BL BLB W_4_29_1 W_4_29_1_bar CIM_cell
X4982 I4292 O_4_29_2_2 WL_4_2 BL BLB W_4_29_2 W_4_29_2_bar CIM_cell
X4983 I4292 O_4_29_2_3 WL_4_2 BL BLB W_4_29_3 W_4_29_3_bar CIM_cell
X4984 I4292 O_4_29_2_4 WL_4_2 BL BLB W_4_29_4 W_4_29_4_bar CIM_cell
X4991 I4293 O_4_29_3_1 WL_4_3 BL BLB W_4_29_1 W_4_29_1_bar CIM_cell
X4992 I4293 O_4_29_3_2 WL_4_3 BL BLB W_4_29_2 W_4_29_2_bar CIM_cell
X4993 I4293 O_4_29_3_3 WL_4_3 BL BLB W_4_29_3 W_4_29_3_bar CIM_cell
X4994 I4293 O_4_29_3_4 WL_4_3 BL BLB W_4_29_4 W_4_29_4_bar CIM_cell
X5001 I4294 O_4_29_4_1 WL_4_4 BL BLB W_4_29_1 W_4_29_1_bar CIM_cell
X5002 I4294 O_4_29_4_2 WL_4_4 BL BLB W_4_29_2 W_4_29_2_bar CIM_cell
X5003 I4294 O_4_29_4_3 WL_4_4 BL BLB W_4_29_3 W_4_29_3_bar CIM_cell
X5004 I4294 O_4_29_4_4 WL_4_4 BL BLB W_4_29_4 W_4_29_4_bar CIM_cell
X5011 I4301 O_4_30_1_1 WL_4_1 BL BLB W_4_30_1 W_4_30_1_bar CIM_cell
X5012 I4301 O_4_30_1_2 WL_4_1 BL BLB W_4_30_2 W_4_30_2_bar CIM_cell
X5013 I4301 O_4_30_1_3 WL_4_1 BL BLB W_4_30_3 W_4_30_3_bar CIM_cell
X5014 I4301 O_4_30_1_4 WL_4_1 BL BLB W_4_30_4 W_4_30_4_bar CIM_cell
X5021 I4302 O_4_30_2_1 WL_4_2 BL BLB W_4_30_1 W_4_30_1_bar CIM_cell
X5022 I4302 O_4_30_2_2 WL_4_2 BL BLB W_4_30_2 W_4_30_2_bar CIM_cell
X5023 I4302 O_4_30_2_3 WL_4_2 BL BLB W_4_30_3 W_4_30_3_bar CIM_cell
X5024 I4302 O_4_30_2_4 WL_4_2 BL BLB W_4_30_4 W_4_30_4_bar CIM_cell
X5031 I4303 O_4_30_3_1 WL_4_3 BL BLB W_4_30_1 W_4_30_1_bar CIM_cell
X5032 I4303 O_4_30_3_2 WL_4_3 BL BLB W_4_30_2 W_4_30_2_bar CIM_cell
X5033 I4303 O_4_30_3_3 WL_4_3 BL BLB W_4_30_3 W_4_30_3_bar CIM_cell
X5034 I4303 O_4_30_3_4 WL_4_3 BL BLB W_4_30_4 W_4_30_4_bar CIM_cell
X5041 I4304 O_4_30_4_1 WL_4_4 BL BLB W_4_30_1 W_4_30_1_bar CIM_cell
X5042 I4304 O_4_30_4_2 WL_4_4 BL BLB W_4_30_2 W_4_30_2_bar CIM_cell
X5043 I4304 O_4_30_4_3 WL_4_4 BL BLB W_4_30_3 W_4_30_3_bar CIM_cell
X5044 I4304 O_4_30_4_4 WL_4_4 BL BLB W_4_30_4 W_4_30_4_bar CIM_cell
X5051 I4311 O_4_31_1_1 WL_4_1 BL BLB W_4_31_1 W_4_31_1_bar CIM_cell
X5052 I4311 O_4_31_1_2 WL_4_1 BL BLB W_4_31_2 W_4_31_2_bar CIM_cell
X5053 I4311 O_4_31_1_3 WL_4_1 BL BLB W_4_31_3 W_4_31_3_bar CIM_cell
X5054 I4311 O_4_31_1_4 WL_4_1 BL BLB W_4_31_4 W_4_31_4_bar CIM_cell
X5061 I4312 O_4_31_2_1 WL_4_2 BL BLB W_4_31_1 W_4_31_1_bar CIM_cell
X5062 I4312 O_4_31_2_2 WL_4_2 BL BLB W_4_31_2 W_4_31_2_bar CIM_cell
X5063 I4312 O_4_31_2_3 WL_4_2 BL BLB W_4_31_3 W_4_31_3_bar CIM_cell
X5064 I4312 O_4_31_2_4 WL_4_2 BL BLB W_4_31_4 W_4_31_4_bar CIM_cell
X5071 I4313 O_4_31_3_1 WL_4_3 BL BLB W_4_31_1 W_4_31_1_bar CIM_cell
X5072 I4313 O_4_31_3_2 WL_4_3 BL BLB W_4_31_2 W_4_31_2_bar CIM_cell
X5073 I4313 O_4_31_3_3 WL_4_3 BL BLB W_4_31_3 W_4_31_3_bar CIM_cell
X5074 I4313 O_4_31_3_4 WL_4_3 BL BLB W_4_31_4 W_4_31_4_bar CIM_cell
X5081 I4314 O_4_31_4_1 WL_4_4 BL BLB W_4_31_1 W_4_31_1_bar CIM_cell
X5082 I4314 O_4_31_4_2 WL_4_4 BL BLB W_4_31_2 W_4_31_2_bar CIM_cell
X5083 I4314 O_4_31_4_3 WL_4_4 BL BLB W_4_31_3 W_4_31_3_bar CIM_cell
X5084 I4314 O_4_31_4_4 WL_4_4 BL BLB W_4_31_4 W_4_31_4_bar CIM_cell
X5091 I4321 O_4_32_1_1 WL_4_1 BL BLB W_4_32_1 W_4_32_1_bar CIM_cell
X5092 I4321 O_4_32_1_2 WL_4_1 BL BLB W_4_32_2 W_4_32_2_bar CIM_cell
X5093 I4321 O_4_32_1_3 WL_4_1 BL BLB W_4_32_3 W_4_32_3_bar CIM_cell
X5094 I4321 O_4_32_1_4 WL_4_1 BL BLB W_4_32_4 W_4_32_4_bar CIM_cell
X5101 I4322 O_4_32_2_1 WL_4_2 BL BLB W_4_32_1 W_4_32_1_bar CIM_cell
X5102 I4322 O_4_32_2_2 WL_4_2 BL BLB W_4_32_2 W_4_32_2_bar CIM_cell
X5103 I4322 O_4_32_2_3 WL_4_2 BL BLB W_4_32_3 W_4_32_3_bar CIM_cell
X5104 I4322 O_4_32_2_4 WL_4_2 BL BLB W_4_32_4 W_4_32_4_bar CIM_cell
X5111 I4323 O_4_32_3_1 WL_4_3 BL BLB W_4_32_1 W_4_32_1_bar CIM_cell
X5112 I4323 O_4_32_3_2 WL_4_3 BL BLB W_4_32_2 W_4_32_2_bar CIM_cell
X5113 I4323 O_4_32_3_3 WL_4_3 BL BLB W_4_32_3 W_4_32_3_bar CIM_cell
X5114 I4323 O_4_32_3_4 WL_4_3 BL BLB W_4_32_4 W_4_32_4_bar CIM_cell
X5121 I4324 O_4_32_4_1 WL_4_4 BL BLB W_4_32_1 W_4_32_1_bar CIM_cell
X5122 I4324 O_4_32_4_2 WL_4_4 BL BLB W_4_32_2 W_4_32_2_bar CIM_cell
X5123 I4324 O_4_32_4_3 WL_4_4 BL BLB W_4_32_3 W_4_32_3_bar CIM_cell
X5124 I4324 O_4_32_4_4 WL_4_4 BL BLB W_4_32_4 W_4_32_4_bar CIM_cell


***-----------------------***
***      sub-circuit      ***
***-----------------------***

* // QB : weight 
* // input 
* // output 
* .subckt CIM_cell Input Output WL BL BLB q qb
*     X01 WL BL BLB q qb SRAM_6T
*     X02 qb Input Output NOR_2
* .ends

.subckt CIM_cell Input Output WL BL BLB q qb
    X01 WL BL BLB q qb SRAM_6T
    X02 q q q1 NOR_2
    X03 Input Input Input1 NOR_2
    X04 q1 Input1 Output NOR_2
.ends


.subckt SRAM_6T WL BL BLB q qb
    MP1 q   qb  VDD VDD pmos_sram m=1
    MP2 qb  q   VDD VDD pmos_sram m=1
    MN1 q   qb  GND GND nmos_sram m=1
    MN2 qb  q   GND GND nmos_sram m=1
    MN3 BL  WL  q   GND nmos_sram m=1
    MN4 qb  WL  BLB GND nmos_sram m=1
.ends

.subckt NOR_2 A B Y
    MP1 N1  A   VDD VDD pmos_lvt m=1
    MP2 Y   B   N1  VDD pmos_lvt m=1
    MN1 Y   A   GND GND nmos_lvt m=1
    MN2 Y   B   GND GND nmos_lvt m=1
.ends

.subckt Buffer in out
    X_INV1 in   in_b INV
    X_INV2 in_b out  INV
.ends

.subckt INV in out
    Mp  out  in  VDD  VDD  pmos_lvt  m=1
    Mn  out  in  GND  GND  nmos_lvt  m=1
.ends

* Example .IC file for initializing SRAM weights
.IC V(W_1_1_1) = 0 V(W_1_1_1_bar) = 1
.IC V(W_1_1_2) = 1 V(W_1_1_2_bar) = 0
.IC V(W_1_1_3) = 0 V(W_1_1_3_bar) = 1
.IC V(W_1_1_4) = 1 V(W_1_1_4_bar) = 0
.IC V(W_1_2_1) = 0 V(W_1_2_1_bar) = 1
.IC V(W_1_2_2) = 1 V(W_1_2_2_bar) = 0
.IC V(W_1_2_3) = 0 V(W_1_2_3_bar) = 1
.IC V(W_1_2_4) = 1 V(W_1_2_4_bar) = 0
.IC V(W_1_3_1) = 0 V(W_1_3_1_bar) = 1
.IC V(W_1_3_2) = 1 V(W_1_3_2_bar) = 0
.IC V(W_1_3_3) = 0 V(W_1_3_3_bar) = 1
.IC V(W_1_3_4) = 1 V(W_1_3_4_bar) = 0
.IC V(W_1_4_1) = 0 V(W_1_4_1_bar) = 1
.IC V(W_1_4_2) = 1 V(W_1_4_2_bar) = 0
.IC V(W_1_4_3) = 0 V(W_1_4_3_bar) = 1
.IC V(W_1_4_4) = 1 V(W_1_4_4_bar) = 0
.IC V(W_1_5_1) = 0 V(W_1_5_1_bar) = 1
.IC V(W_1_5_2) = 1 V(W_1_5_2_bar) = 0
.IC V(W_1_5_3) = 0 V(W_1_5_3_bar) = 1
.IC V(W_1_5_4) = 1 V(W_1_5_4_bar) = 0
.IC V(W_1_6_1) = 0 V(W_1_6_1_bar) = 1
.IC V(W_1_6_2) = 1 V(W_1_6_2_bar) = 0
.IC V(W_1_6_3) = 0 V(W_1_6_3_bar) = 1
.IC V(W_1_6_4) = 1 V(W_1_6_4_bar) = 0
.IC V(W_1_7_1) = 0 V(W_1_7_1_bar) = 1
.IC V(W_1_7_2) = 1 V(W_1_7_2_bar) = 0
.IC V(W_1_7_3) = 0 V(W_1_7_3_bar) = 1
.IC V(W_1_7_4) = 1 V(W_1_7_4_bar) = 0
.IC V(W_1_8_1) = 0 V(W_1_8_1_bar) = 1
.IC V(W_1_8_2) = 1 V(W_1_8_2_bar) = 0
.IC V(W_1_8_3) = 0 V(W_1_8_3_bar) = 1
.IC V(W_1_8_4) = 1 V(W_1_8_4_bar) = 0
.IC V(W_1_9_1) = 0 V(W_1_9_1_bar) = 1
.IC V(W_1_9_2) = 1 V(W_1_9_2_bar) = 0
.IC V(W_1_9_3) = 0 V(W_1_9_3_bar) = 1
.IC V(W_1_9_4) = 1 V(W_1_9_4_bar) = 0
.IC V(W_1_10_1) = 0 V(W_1_10_1_bar) = 1
.IC V(W_1_10_2) = 1 V(W_1_10_2_bar) = 0
.IC V(W_1_10_3) = 0 V(W_1_10_3_bar) = 1
.IC V(W_1_10_4) = 1 V(W_1_10_4_bar) = 0
.IC V(W_1_11_1) = 0 V(W_1_11_1_bar) = 1
.IC V(W_1_11_2) = 1 V(W_1_11_2_bar) = 0
.IC V(W_1_11_3) = 0 V(W_1_11_3_bar) = 1
.IC V(W_1_11_4) = 1 V(W_1_11_4_bar) = 0
.IC V(W_1_12_1) = 0 V(W_1_12_1_bar) = 1
.IC V(W_1_12_2) = 1 V(W_1_12_2_bar) = 0
.IC V(W_1_12_3) = 0 V(W_1_12_3_bar) = 1
.IC V(W_1_12_4) = 1 V(W_1_12_4_bar) = 0
.IC V(W_1_13_1) = 0 V(W_1_13_1_bar) = 1
.IC V(W_1_13_2) = 1 V(W_1_13_2_bar) = 0
.IC V(W_1_13_3) = 0 V(W_1_13_3_bar) = 1
.IC V(W_1_13_4) = 1 V(W_1_13_4_bar) = 0
.IC V(W_1_14_1) = 0 V(W_1_14_1_bar) = 1
.IC V(W_1_14_2) = 1 V(W_1_14_2_bar) = 0
.IC V(W_1_14_3) = 0 V(W_1_14_3_bar) = 1
.IC V(W_1_14_4) = 1 V(W_1_14_4_bar) = 0
.IC V(W_1_15_1) = 0 V(W_1_15_1_bar) = 1
.IC V(W_1_15_2) = 1 V(W_1_15_2_bar) = 0
.IC V(W_1_15_3) = 0 V(W_1_15_3_bar) = 1
.IC V(W_1_15_4) = 1 V(W_1_15_4_bar) = 0
.IC V(W_1_16_1) = 0 V(W_1_16_1_bar) = 1
.IC V(W_1_16_2) = 1 V(W_1_16_2_bar) = 0
.IC V(W_1_16_3) = 0 V(W_1_16_3_bar) = 1
.IC V(W_1_16_4) = 1 V(W_1_16_4_bar) = 0
.IC V(W_1_17_1) = 0 V(W_1_17_1_bar) = 1
.IC V(W_1_17_2) = 1 V(W_1_17_2_bar) = 0
.IC V(W_1_17_3) = 0 V(W_1_17_3_bar) = 1
.IC V(W_1_17_4) = 1 V(W_1_17_4_bar) = 0
.IC V(W_1_18_1) = 0 V(W_1_18_1_bar) = 1
.IC V(W_1_18_2) = 1 V(W_1_18_2_bar) = 0
.IC V(W_1_18_3) = 0 V(W_1_18_3_bar) = 1
.IC V(W_1_18_4) = 1 V(W_1_18_4_bar) = 0
.IC V(W_1_19_1) = 0 V(W_1_19_1_bar) = 1
.IC V(W_1_19_2) = 1 V(W_1_19_2_bar) = 0
.IC V(W_1_19_3) = 0 V(W_1_19_3_bar) = 1
.IC V(W_1_19_4) = 1 V(W_1_19_4_bar) = 0
.IC V(W_1_20_1) = 0 V(W_1_20_1_bar) = 1
.IC V(W_1_20_2) = 1 V(W_1_20_2_bar) = 0
.IC V(W_1_20_3) = 0 V(W_1_20_3_bar) = 1
.IC V(W_1_20_4) = 1 V(W_1_20_4_bar) = 0
.IC V(W_1_21_1) = 0 V(W_1_21_1_bar) = 1
.IC V(W_1_21_2) = 1 V(W_1_21_2_bar) = 0
.IC V(W_1_21_3) = 0 V(W_1_21_3_bar) = 1
.IC V(W_1_21_4) = 1 V(W_1_21_4_bar) = 0
.IC V(W_1_22_1) = 0 V(W_1_22_1_bar) = 1
.IC V(W_1_22_2) = 1 V(W_1_22_2_bar) = 0
.IC V(W_1_22_3) = 0 V(W_1_22_3_bar) = 1
.IC V(W_1_22_4) = 1 V(W_1_22_4_bar) = 0
.IC V(W_1_23_1) = 0 V(W_1_23_1_bar) = 1
.IC V(W_1_23_2) = 1 V(W_1_23_2_bar) = 0
.IC V(W_1_23_3) = 0 V(W_1_23_3_bar) = 1
.IC V(W_1_23_4) = 1 V(W_1_23_4_bar) = 0
.IC V(W_1_24_1) = 0 V(W_1_24_1_bar) = 1
.IC V(W_1_24_2) = 1 V(W_1_24_2_bar) = 0
.IC V(W_1_24_3) = 0 V(W_1_24_3_bar) = 1
.IC V(W_1_24_4) = 1 V(W_1_24_4_bar) = 0
.IC V(W_1_25_1) = 0 V(W_1_25_1_bar) = 1
.IC V(W_1_25_2) = 1 V(W_1_25_2_bar) = 0
.IC V(W_1_25_3) = 0 V(W_1_25_3_bar) = 1
.IC V(W_1_25_4) = 1 V(W_1_25_4_bar) = 0
.IC V(W_1_26_1) = 0 V(W_1_26_1_bar) = 1
.IC V(W_1_26_2) = 1 V(W_1_26_2_bar) = 0
.IC V(W_1_26_3) = 0 V(W_1_26_3_bar) = 1
.IC V(W_1_26_4) = 1 V(W_1_26_4_bar) = 0
.IC V(W_1_27_1) = 0 V(W_1_27_1_bar) = 1
.IC V(W_1_27_2) = 1 V(W_1_27_2_bar) = 0
.IC V(W_1_27_3) = 0 V(W_1_27_3_bar) = 1
.IC V(W_1_27_4) = 1 V(W_1_27_4_bar) = 0
.IC V(W_1_28_1) = 0 V(W_1_28_1_bar) = 1
.IC V(W_1_28_2) = 1 V(W_1_28_2_bar) = 0
.IC V(W_1_28_3) = 0 V(W_1_28_3_bar) = 1
.IC V(W_1_28_4) = 1 V(W_1_28_4_bar) = 0
.IC V(W_1_29_1) = 0 V(W_1_29_1_bar) = 1
.IC V(W_1_29_2) = 1 V(W_1_29_2_bar) = 0
.IC V(W_1_29_3) = 0 V(W_1_29_3_bar) = 1
.IC V(W_1_29_4) = 1 V(W_1_29_4_bar) = 0
.IC V(W_1_30_1) = 0 V(W_1_30_1_bar) = 1
.IC V(W_1_30_2) = 1 V(W_1_30_2_bar) = 0
.IC V(W_1_30_3) = 0 V(W_1_30_3_bar) = 1
.IC V(W_1_30_4) = 1 V(W_1_30_4_bar) = 0
.IC V(W_1_31_1) = 0 V(W_1_31_1_bar) = 1
.IC V(W_1_31_2) = 1 V(W_1_31_2_bar) = 0
.IC V(W_1_31_3) = 0 V(W_1_31_3_bar) = 1
.IC V(W_1_31_4) = 1 V(W_1_31_4_bar) = 0
.IC V(W_1_32_1) = 0 V(W_1_32_1_bar) = 1
.IC V(W_1_32_2) = 1 V(W_1_32_2_bar) = 0
.IC V(W_1_32_3) = 0 V(W_1_32_3_bar) = 1
.IC V(W_1_32_4) = 1 V(W_1_32_4_bar) = 0
.IC V(W_2_1_1) = 0 V(W_2_1_1_bar) = 1
.IC V(W_2_1_2) = 1 V(W_2_1_2_bar) = 0
.IC V(W_2_1_3) = 0 V(W_2_1_3_bar) = 1
.IC V(W_2_1_4) = 1 V(W_2_1_4_bar) = 0
.IC V(W_2_2_1) = 0 V(W_2_2_1_bar) = 1
.IC V(W_2_2_2) = 1 V(W_2_2_2_bar) = 0
.IC V(W_2_2_3) = 0 V(W_2_2_3_bar) = 1
.IC V(W_2_2_4) = 1 V(W_2_2_4_bar) = 0
.IC V(W_2_3_1) = 0 V(W_2_3_1_bar) = 1
.IC V(W_2_3_2) = 1 V(W_2_3_2_bar) = 0
.IC V(W_2_3_3) = 0 V(W_2_3_3_bar) = 1
.IC V(W_2_3_4) = 1 V(W_2_3_4_bar) = 0
.IC V(W_2_4_1) = 0 V(W_2_4_1_bar) = 1
.IC V(W_2_4_2) = 1 V(W_2_4_2_bar) = 0
.IC V(W_2_4_3) = 0 V(W_2_4_3_bar) = 1
.IC V(W_2_4_4) = 1 V(W_2_4_4_bar) = 0
.IC V(W_2_5_1) = 0 V(W_2_5_1_bar) = 1
.IC V(W_2_5_2) = 1 V(W_2_5_2_bar) = 0
.IC V(W_2_5_3) = 0 V(W_2_5_3_bar) = 1
.IC V(W_2_5_4) = 1 V(W_2_5_4_bar) = 0
.IC V(W_2_6_1) = 0 V(W_2_6_1_bar) = 1
.IC V(W_2_6_2) = 1 V(W_2_6_2_bar) = 0
.IC V(W_2_6_3) = 0 V(W_2_6_3_bar) = 1
.IC V(W_2_6_4) = 1 V(W_2_6_4_bar) = 0
.IC V(W_2_7_1) = 0 V(W_2_7_1_bar) = 1
.IC V(W_2_7_2) = 1 V(W_2_7_2_bar) = 0
.IC V(W_2_7_3) = 0 V(W_2_7_3_bar) = 1
.IC V(W_2_7_4) = 1 V(W_2_7_4_bar) = 0
.IC V(W_2_8_1) = 0 V(W_2_8_1_bar) = 1
.IC V(W_2_8_2) = 1 V(W_2_8_2_bar) = 0
.IC V(W_2_8_3) = 0 V(W_2_8_3_bar) = 1
.IC V(W_2_8_4) = 1 V(W_2_8_4_bar) = 0
.IC V(W_2_9_1) = 0 V(W_2_9_1_bar) = 1
.IC V(W_2_9_2) = 1 V(W_2_9_2_bar) = 0
.IC V(W_2_9_3) = 0 V(W_2_9_3_bar) = 1
.IC V(W_2_9_4) = 1 V(W_2_9_4_bar) = 0
.IC V(W_2_10_1) = 0 V(W_2_10_1_bar) = 1
.IC V(W_2_10_2) = 1 V(W_2_10_2_bar) = 0
.IC V(W_2_10_3) = 0 V(W_2_10_3_bar) = 1
.IC V(W_2_10_4) = 1 V(W_2_10_4_bar) = 0
.IC V(W_2_11_1) = 0 V(W_2_11_1_bar) = 1
.IC V(W_2_11_2) = 1 V(W_2_11_2_bar) = 0
.IC V(W_2_11_3) = 0 V(W_2_11_3_bar) = 1
.IC V(W_2_11_4) = 1 V(W_2_11_4_bar) = 0
.IC V(W_2_12_1) = 0 V(W_2_12_1_bar) = 1
.IC V(W_2_12_2) = 1 V(W_2_12_2_bar) = 0
.IC V(W_2_12_3) = 0 V(W_2_12_3_bar) = 1
.IC V(W_2_12_4) = 1 V(W_2_12_4_bar) = 0
.IC V(W_2_13_1) = 0 V(W_2_13_1_bar) = 1
.IC V(W_2_13_2) = 1 V(W_2_13_2_bar) = 0
.IC V(W_2_13_3) = 0 V(W_2_13_3_bar) = 1
.IC V(W_2_13_4) = 1 V(W_2_13_4_bar) = 0
.IC V(W_2_14_1) = 0 V(W_2_14_1_bar) = 1
.IC V(W_2_14_2) = 1 V(W_2_14_2_bar) = 0
.IC V(W_2_14_3) = 0 V(W_2_14_3_bar) = 1
.IC V(W_2_14_4) = 1 V(W_2_14_4_bar) = 0
.IC V(W_2_15_1) = 0 V(W_2_15_1_bar) = 1
.IC V(W_2_15_2) = 1 V(W_2_15_2_bar) = 0
.IC V(W_2_15_3) = 0 V(W_2_15_3_bar) = 1
.IC V(W_2_15_4) = 1 V(W_2_15_4_bar) = 0
.IC V(W_2_16_1) = 0 V(W_2_16_1_bar) = 1
.IC V(W_2_16_2) = 1 V(W_2_16_2_bar) = 0
.IC V(W_2_16_3) = 0 V(W_2_16_3_bar) = 1
.IC V(W_2_16_4) = 1 V(W_2_16_4_bar) = 0
.IC V(W_2_17_1) = 0 V(W_2_17_1_bar) = 1
.IC V(W_2_17_2) = 1 V(W_2_17_2_bar) = 0
.IC V(W_2_17_3) = 0 V(W_2_17_3_bar) = 1
.IC V(W_2_17_4) = 1 V(W_2_17_4_bar) = 0
.IC V(W_2_18_1) = 0 V(W_2_18_1_bar) = 1
.IC V(W_2_18_2) = 1 V(W_2_18_2_bar) = 0
.IC V(W_2_18_3) = 0 V(W_2_18_3_bar) = 1
.IC V(W_2_18_4) = 1 V(W_2_18_4_bar) = 0
.IC V(W_2_19_1) = 0 V(W_2_19_1_bar) = 1
.IC V(W_2_19_2) = 1 V(W_2_19_2_bar) = 0
.IC V(W_2_19_3) = 0 V(W_2_19_3_bar) = 1
.IC V(W_2_19_4) = 1 V(W_2_19_4_bar) = 0
.IC V(W_2_20_1) = 0 V(W_2_20_1_bar) = 1
.IC V(W_2_20_2) = 1 V(W_2_20_2_bar) = 0
.IC V(W_2_20_3) = 0 V(W_2_20_3_bar) = 1
.IC V(W_2_20_4) = 1 V(W_2_20_4_bar) = 0
.IC V(W_2_21_1) = 0 V(W_2_21_1_bar) = 1
.IC V(W_2_21_2) = 1 V(W_2_21_2_bar) = 0
.IC V(W_2_21_3) = 0 V(W_2_21_3_bar) = 1
.IC V(W_2_21_4) = 1 V(W_2_21_4_bar) = 0
.IC V(W_2_22_1) = 0 V(W_2_22_1_bar) = 1
.IC V(W_2_22_2) = 1 V(W_2_22_2_bar) = 0
.IC V(W_2_22_3) = 0 V(W_2_22_3_bar) = 1
.IC V(W_2_22_4) = 1 V(W_2_22_4_bar) = 0
.IC V(W_2_23_1) = 0 V(W_2_23_1_bar) = 1
.IC V(W_2_23_2) = 1 V(W_2_23_2_bar) = 0
.IC V(W_2_23_3) = 0 V(W_2_23_3_bar) = 1
.IC V(W_2_23_4) = 1 V(W_2_23_4_bar) = 0
.IC V(W_2_24_1) = 0 V(W_2_24_1_bar) = 1
.IC V(W_2_24_2) = 1 V(W_2_24_2_bar) = 0
.IC V(W_2_24_3) = 0 V(W_2_24_3_bar) = 1
.IC V(W_2_24_4) = 1 V(W_2_24_4_bar) = 0
.IC V(W_2_25_1) = 0 V(W_2_25_1_bar) = 1
.IC V(W_2_25_2) = 1 V(W_2_25_2_bar) = 0
.IC V(W_2_25_3) = 0 V(W_2_25_3_bar) = 1
.IC V(W_2_25_4) = 1 V(W_2_25_4_bar) = 0
.IC V(W_2_26_1) = 0 V(W_2_26_1_bar) = 1
.IC V(W_2_26_2) = 1 V(W_2_26_2_bar) = 0
.IC V(W_2_26_3) = 0 V(W_2_26_3_bar) = 1
.IC V(W_2_26_4) = 1 V(W_2_26_4_bar) = 0
.IC V(W_2_27_1) = 0 V(W_2_27_1_bar) = 1
.IC V(W_2_27_2) = 1 V(W_2_27_2_bar) = 0
.IC V(W_2_27_3) = 0 V(W_2_27_3_bar) = 1
.IC V(W_2_27_4) = 1 V(W_2_27_4_bar) = 0
.IC V(W_2_28_1) = 0 V(W_2_28_1_bar) = 1
.IC V(W_2_28_2) = 1 V(W_2_28_2_bar) = 0
.IC V(W_2_28_3) = 0 V(W_2_28_3_bar) = 1
.IC V(W_2_28_4) = 1 V(W_2_28_4_bar) = 0
.IC V(W_2_29_1) = 0 V(W_2_29_1_bar) = 1
.IC V(W_2_29_2) = 1 V(W_2_29_2_bar) = 0
.IC V(W_2_29_3) = 0 V(W_2_29_3_bar) = 1
.IC V(W_2_29_4) = 1 V(W_2_29_4_bar) = 0
.IC V(W_2_30_1) = 0 V(W_2_30_1_bar) = 1
.IC V(W_2_30_2) = 1 V(W_2_30_2_bar) = 0
.IC V(W_2_30_3) = 0 V(W_2_30_3_bar) = 1
.IC V(W_2_30_4) = 1 V(W_2_30_4_bar) = 0
.IC V(W_2_31_1) = 0 V(W_2_31_1_bar) = 1
.IC V(W_2_31_2) = 1 V(W_2_31_2_bar) = 0
.IC V(W_2_31_3) = 0 V(W_2_31_3_bar) = 1
.IC V(W_2_31_4) = 1 V(W_2_31_4_bar) = 0
.IC V(W_2_32_1) = 0 V(W_2_32_1_bar) = 1
.IC V(W_2_32_2) = 1 V(W_2_32_2_bar) = 0
.IC V(W_2_32_3) = 0 V(W_2_32_3_bar) = 1
.IC V(W_2_32_4) = 1 V(W_2_32_4_bar) = 0
.IC V(W_3_1_1) = 0 V(W_3_1_1_bar) = 1
.IC V(W_3_1_2) = 1 V(W_3_1_2_bar) = 0
.IC V(W_3_1_3) = 0 V(W_3_1_3_bar) = 1
.IC V(W_3_1_4) = 1 V(W_3_1_4_bar) = 0
.IC V(W_3_2_1) = 0 V(W_3_2_1_bar) = 1
.IC V(W_3_2_2) = 1 V(W_3_2_2_bar) = 0
.IC V(W_3_2_3) = 0 V(W_3_2_3_bar) = 1
.IC V(W_3_2_4) = 1 V(W_3_2_4_bar) = 0
.IC V(W_3_3_1) = 0 V(W_3_3_1_bar) = 1
.IC V(W_3_3_2) = 1 V(W_3_3_2_bar) = 0
.IC V(W_3_3_3) = 0 V(W_3_3_3_bar) = 1
.IC V(W_3_3_4) = 1 V(W_3_3_4_bar) = 0
.IC V(W_3_4_1) = 0 V(W_3_4_1_bar) = 1
.IC V(W_3_4_2) = 1 V(W_3_4_2_bar) = 0
.IC V(W_3_4_3) = 0 V(W_3_4_3_bar) = 1
.IC V(W_3_4_4) = 1 V(W_3_4_4_bar) = 0
.IC V(W_3_5_1) = 0 V(W_3_5_1_bar) = 1
.IC V(W_3_5_2) = 1 V(W_3_5_2_bar) = 0
.IC V(W_3_5_3) = 0 V(W_3_5_3_bar) = 1
.IC V(W_3_5_4) = 1 V(W_3_5_4_bar) = 0
.IC V(W_3_6_1) = 0 V(W_3_6_1_bar) = 1
.IC V(W_3_6_2) = 1 V(W_3_6_2_bar) = 0
.IC V(W_3_6_3) = 0 V(W_3_6_3_bar) = 1
.IC V(W_3_6_4) = 1 V(W_3_6_4_bar) = 0
.IC V(W_3_7_1) = 0 V(W_3_7_1_bar) = 1
.IC V(W_3_7_2) = 1 V(W_3_7_2_bar) = 0
.IC V(W_3_7_3) = 0 V(W_3_7_3_bar) = 1
.IC V(W_3_7_4) = 1 V(W_3_7_4_bar) = 0
.IC V(W_3_8_1) = 0 V(W_3_8_1_bar) = 1
.IC V(W_3_8_2) = 1 V(W_3_8_2_bar) = 0
.IC V(W_3_8_3) = 0 V(W_3_8_3_bar) = 1
.IC V(W_3_8_4) = 1 V(W_3_8_4_bar) = 0
.IC V(W_3_9_1) = 0 V(W_3_9_1_bar) = 1
.IC V(W_3_9_2) = 1 V(W_3_9_2_bar) = 0
.IC V(W_3_9_3) = 0 V(W_3_9_3_bar) = 1
.IC V(W_3_9_4) = 1 V(W_3_9_4_bar) = 0
.IC V(W_3_10_1) = 0 V(W_3_10_1_bar) = 1
.IC V(W_3_10_2) = 1 V(W_3_10_2_bar) = 0
.IC V(W_3_10_3) = 0 V(W_3_10_3_bar) = 1
.IC V(W_3_10_4) = 1 V(W_3_10_4_bar) = 0
.IC V(W_3_11_1) = 0 V(W_3_11_1_bar) = 1
.IC V(W_3_11_2) = 1 V(W_3_11_2_bar) = 0
.IC V(W_3_11_3) = 0 V(W_3_11_3_bar) = 1
.IC V(W_3_11_4) = 1 V(W_3_11_4_bar) = 0
.IC V(W_3_12_1) = 0 V(W_3_12_1_bar) = 1
.IC V(W_3_12_2) = 1 V(W_3_12_2_bar) = 0
.IC V(W_3_12_3) = 0 V(W_3_12_3_bar) = 1
.IC V(W_3_12_4) = 1 V(W_3_12_4_bar) = 0
.IC V(W_3_13_1) = 0 V(W_3_13_1_bar) = 1
.IC V(W_3_13_2) = 1 V(W_3_13_2_bar) = 0
.IC V(W_3_13_3) = 0 V(W_3_13_3_bar) = 1
.IC V(W_3_13_4) = 1 V(W_3_13_4_bar) = 0
.IC V(W_3_14_1) = 0 V(W_3_14_1_bar) = 1
.IC V(W_3_14_2) = 1 V(W_3_14_2_bar) = 0
.IC V(W_3_14_3) = 0 V(W_3_14_3_bar) = 1
.IC V(W_3_14_4) = 1 V(W_3_14_4_bar) = 0
.IC V(W_3_15_1) = 0 V(W_3_15_1_bar) = 1
.IC V(W_3_15_2) = 1 V(W_3_15_2_bar) = 0
.IC V(W_3_15_3) = 0 V(W_3_15_3_bar) = 1
.IC V(W_3_15_4) = 1 V(W_3_15_4_bar) = 0
.IC V(W_3_16_1) = 0 V(W_3_16_1_bar) = 1
.IC V(W_3_16_2) = 1 V(W_3_16_2_bar) = 0
.IC V(W_3_16_3) = 0 V(W_3_16_3_bar) = 1
.IC V(W_3_16_4) = 1 V(W_3_16_4_bar) = 0
.IC V(W_3_17_1) = 0 V(W_3_17_1_bar) = 1
.IC V(W_3_17_2) = 1 V(W_3_17_2_bar) = 0
.IC V(W_3_17_3) = 0 V(W_3_17_3_bar) = 1
.IC V(W_3_17_4) = 1 V(W_3_17_4_bar) = 0
.IC V(W_3_18_1) = 0 V(W_3_18_1_bar) = 1
.IC V(W_3_18_2) = 1 V(W_3_18_2_bar) = 0
.IC V(W_3_18_3) = 0 V(W_3_18_3_bar) = 1
.IC V(W_3_18_4) = 1 V(W_3_18_4_bar) = 0
.IC V(W_3_19_1) = 0 V(W_3_19_1_bar) = 1
.IC V(W_3_19_2) = 1 V(W_3_19_2_bar) = 0
.IC V(W_3_19_3) = 0 V(W_3_19_3_bar) = 1
.IC V(W_3_19_4) = 1 V(W_3_19_4_bar) = 0
.IC V(W_3_20_1) = 0 V(W_3_20_1_bar) = 1
.IC V(W_3_20_2) = 1 V(W_3_20_2_bar) = 0
.IC V(W_3_20_3) = 0 V(W_3_20_3_bar) = 1
.IC V(W_3_20_4) = 1 V(W_3_20_4_bar) = 0
.IC V(W_3_21_1) = 0 V(W_3_21_1_bar) = 1
.IC V(W_3_21_2) = 1 V(W_3_21_2_bar) = 0
.IC V(W_3_21_3) = 0 V(W_3_21_3_bar) = 1
.IC V(W_3_21_4) = 1 V(W_3_21_4_bar) = 0
.IC V(W_3_22_1) = 0 V(W_3_22_1_bar) = 1
.IC V(W_3_22_2) = 1 V(W_3_22_2_bar) = 0
.IC V(W_3_22_3) = 0 V(W_3_22_3_bar) = 1
.IC V(W_3_22_4) = 1 V(W_3_22_4_bar) = 0
.IC V(W_3_23_1) = 0 V(W_3_23_1_bar) = 1
.IC V(W_3_23_2) = 1 V(W_3_23_2_bar) = 0
.IC V(W_3_23_3) = 0 V(W_3_23_3_bar) = 1
.IC V(W_3_23_4) = 1 V(W_3_23_4_bar) = 0
.IC V(W_3_24_1) = 0 V(W_3_24_1_bar) = 1
.IC V(W_3_24_2) = 1 V(W_3_24_2_bar) = 0
.IC V(W_3_24_3) = 0 V(W_3_24_3_bar) = 1
.IC V(W_3_24_4) = 1 V(W_3_24_4_bar) = 0
.IC V(W_3_25_1) = 0 V(W_3_25_1_bar) = 1
.IC V(W_3_25_2) = 1 V(W_3_25_2_bar) = 0
.IC V(W_3_25_3) = 0 V(W_3_25_3_bar) = 1
.IC V(W_3_25_4) = 1 V(W_3_25_4_bar) = 0
.IC V(W_3_26_1) = 0 V(W_3_26_1_bar) = 1
.IC V(W_3_26_2) = 1 V(W_3_26_2_bar) = 0
.IC V(W_3_26_3) = 0 V(W_3_26_3_bar) = 1
.IC V(W_3_26_4) = 1 V(W_3_26_4_bar) = 0
.IC V(W_3_27_1) = 0 V(W_3_27_1_bar) = 1
.IC V(W_3_27_2) = 1 V(W_3_27_2_bar) = 0
.IC V(W_3_27_3) = 0 V(W_3_27_3_bar) = 1
.IC V(W_3_27_4) = 1 V(W_3_27_4_bar) = 0
.IC V(W_3_28_1) = 0 V(W_3_28_1_bar) = 1
.IC V(W_3_28_2) = 1 V(W_3_28_2_bar) = 0
.IC V(W_3_28_3) = 0 V(W_3_28_3_bar) = 1
.IC V(W_3_28_4) = 1 V(W_3_28_4_bar) = 0
.IC V(W_3_29_1) = 0 V(W_3_29_1_bar) = 1
.IC V(W_3_29_2) = 1 V(W_3_29_2_bar) = 0
.IC V(W_3_29_3) = 0 V(W_3_29_3_bar) = 1
.IC V(W_3_29_4) = 1 V(W_3_29_4_bar) = 0
.IC V(W_3_30_1) = 0 V(W_3_30_1_bar) = 1
.IC V(W_3_30_2) = 1 V(W_3_30_2_bar) = 0
.IC V(W_3_30_3) = 0 V(W_3_30_3_bar) = 1
.IC V(W_3_30_4) = 1 V(W_3_30_4_bar) = 0
.IC V(W_3_31_1) = 0 V(W_3_31_1_bar) = 1
.IC V(W_3_31_2) = 1 V(W_3_31_2_bar) = 0
.IC V(W_3_31_3) = 0 V(W_3_31_3_bar) = 1
.IC V(W_3_31_4) = 1 V(W_3_31_4_bar) = 0
.IC V(W_3_32_1) = 0 V(W_3_32_1_bar) = 1
.IC V(W_3_32_2) = 1 V(W_3_32_2_bar) = 0
.IC V(W_3_32_3) = 0 V(W_3_32_3_bar) = 1
.IC V(W_3_32_4) = 1 V(W_3_32_4_bar) = 0
.IC V(W_4_1_1) = 0 V(W_4_1_1_bar) = 1
.IC V(W_4_1_2) = 1 V(W_4_1_2_bar) = 0
.IC V(W_4_1_3) = 0 V(W_4_1_3_bar) = 1
.IC V(W_4_1_4) = 1 V(W_4_1_4_bar) = 0
.IC V(W_4_2_1) = 0 V(W_4_2_1_bar) = 1
.IC V(W_4_2_2) = 1 V(W_4_2_2_bar) = 0
.IC V(W_4_2_3) = 0 V(W_4_2_3_bar) = 1
.IC V(W_4_2_4) = 1 V(W_4_2_4_bar) = 0
.IC V(W_4_3_1) = 0 V(W_4_3_1_bar) = 1
.IC V(W_4_3_2) = 1 V(W_4_3_2_bar) = 0
.IC V(W_4_3_3) = 0 V(W_4_3_3_bar) = 1
.IC V(W_4_3_4) = 1 V(W_4_3_4_bar) = 0
.IC V(W_4_4_1) = 0 V(W_4_4_1_bar) = 1
.IC V(W_4_4_2) = 1 V(W_4_4_2_bar) = 0
.IC V(W_4_4_3) = 0 V(W_4_4_3_bar) = 1
.IC V(W_4_4_4) = 1 V(W_4_4_4_bar) = 0
.IC V(W_4_5_1) = 0 V(W_4_5_1_bar) = 1
.IC V(W_4_5_2) = 1 V(W_4_5_2_bar) = 0
.IC V(W_4_5_3) = 0 V(W_4_5_3_bar) = 1
.IC V(W_4_5_4) = 1 V(W_4_5_4_bar) = 0
.IC V(W_4_6_1) = 0 V(W_4_6_1_bar) = 1
.IC V(W_4_6_2) = 1 V(W_4_6_2_bar) = 0
.IC V(W_4_6_3) = 0 V(W_4_6_3_bar) = 1
.IC V(W_4_6_4) = 1 V(W_4_6_4_bar) = 0
.IC V(W_4_7_1) = 0 V(W_4_7_1_bar) = 1
.IC V(W_4_7_2) = 1 V(W_4_7_2_bar) = 0
.IC V(W_4_7_3) = 0 V(W_4_7_3_bar) = 1
.IC V(W_4_7_4) = 1 V(W_4_7_4_bar) = 0
.IC V(W_4_8_1) = 0 V(W_4_8_1_bar) = 1
.IC V(W_4_8_2) = 1 V(W_4_8_2_bar) = 0
.IC V(W_4_8_3) = 0 V(W_4_8_3_bar) = 1
.IC V(W_4_8_4) = 1 V(W_4_8_4_bar) = 0
.IC V(W_4_9_1) = 0 V(W_4_9_1_bar) = 1
.IC V(W_4_9_2) = 1 V(W_4_9_2_bar) = 0
.IC V(W_4_9_3) = 0 V(W_4_9_3_bar) = 1
.IC V(W_4_9_4) = 1 V(W_4_9_4_bar) = 0
.IC V(W_4_10_1) = 0 V(W_4_10_1_bar) = 1
.IC V(W_4_10_2) = 1 V(W_4_10_2_bar) = 0
.IC V(W_4_10_3) = 0 V(W_4_10_3_bar) = 1
.IC V(W_4_10_4) = 1 V(W_4_10_4_bar) = 0
.IC V(W_4_11_1) = 0 V(W_4_11_1_bar) = 1
.IC V(W_4_11_2) = 1 V(W_4_11_2_bar) = 0
.IC V(W_4_11_3) = 0 V(W_4_11_3_bar) = 1
.IC V(W_4_11_4) = 1 V(W_4_11_4_bar) = 0
.IC V(W_4_12_1) = 0 V(W_4_12_1_bar) = 1
.IC V(W_4_12_2) = 1 V(W_4_12_2_bar) = 0
.IC V(W_4_12_3) = 0 V(W_4_12_3_bar) = 1
.IC V(W_4_12_4) = 1 V(W_4_12_4_bar) = 0
.IC V(W_4_13_1) = 0 V(W_4_13_1_bar) = 1
.IC V(W_4_13_2) = 1 V(W_4_13_2_bar) = 0
.IC V(W_4_13_3) = 0 V(W_4_13_3_bar) = 1
.IC V(W_4_13_4) = 1 V(W_4_13_4_bar) = 0
.IC V(W_4_14_1) = 0 V(W_4_14_1_bar) = 1
.IC V(W_4_14_2) = 1 V(W_4_14_2_bar) = 0
.IC V(W_4_14_3) = 0 V(W_4_14_3_bar) = 1
.IC V(W_4_14_4) = 1 V(W_4_14_4_bar) = 0
.IC V(W_4_15_1) = 0 V(W_4_15_1_bar) = 1
.IC V(W_4_15_2) = 1 V(W_4_15_2_bar) = 0
.IC V(W_4_15_3) = 0 V(W_4_15_3_bar) = 1
.IC V(W_4_15_4) = 1 V(W_4_15_4_bar) = 0
.IC V(W_4_16_1) = 0 V(W_4_16_1_bar) = 1
.IC V(W_4_16_2) = 1 V(W_4_16_2_bar) = 0
.IC V(W_4_16_3) = 0 V(W_4_16_3_bar) = 1
.IC V(W_4_16_4) = 1 V(W_4_16_4_bar) = 0
.IC V(W_4_17_1) = 0 V(W_4_17_1_bar) = 1
.IC V(W_4_17_2) = 1 V(W_4_17_2_bar) = 0
.IC V(W_4_17_3) = 0 V(W_4_17_3_bar) = 1
.IC V(W_4_17_4) = 1 V(W_4_17_4_bar) = 0
.IC V(W_4_18_1) = 0 V(W_4_18_1_bar) = 1
.IC V(W_4_18_2) = 1 V(W_4_18_2_bar) = 0
.IC V(W_4_18_3) = 0 V(W_4_18_3_bar) = 1
.IC V(W_4_18_4) = 1 V(W_4_18_4_bar) = 0
.IC V(W_4_19_1) = 0 V(W_4_19_1_bar) = 1
.IC V(W_4_19_2) = 1 V(W_4_19_2_bar) = 0
.IC V(W_4_19_3) = 0 V(W_4_19_3_bar) = 1
.IC V(W_4_19_4) = 1 V(W_4_19_4_bar) = 0
.IC V(W_4_20_1) = 0 V(W_4_20_1_bar) = 1
.IC V(W_4_20_2) = 1 V(W_4_20_2_bar) = 0
.IC V(W_4_20_3) = 0 V(W_4_20_3_bar) = 1
.IC V(W_4_20_4) = 1 V(W_4_20_4_bar) = 0
.IC V(W_4_21_1) = 0 V(W_4_21_1_bar) = 1
.IC V(W_4_21_2) = 1 V(W_4_21_2_bar) = 0
.IC V(W_4_21_3) = 0 V(W_4_21_3_bar) = 1
.IC V(W_4_21_4) = 1 V(W_4_21_4_bar) = 0
.IC V(W_4_22_1) = 0 V(W_4_22_1_bar) = 1
.IC V(W_4_22_2) = 1 V(W_4_22_2_bar) = 0
.IC V(W_4_22_3) = 0 V(W_4_22_3_bar) = 1
.IC V(W_4_22_4) = 1 V(W_4_22_4_bar) = 0
.IC V(W_4_23_1) = 0 V(W_4_23_1_bar) = 1
.IC V(W_4_23_2) = 1 V(W_4_23_2_bar) = 0
.IC V(W_4_23_3) = 0 V(W_4_23_3_bar) = 1
.IC V(W_4_23_4) = 1 V(W_4_23_4_bar) = 0
.IC V(W_4_24_1) = 0 V(W_4_24_1_bar) = 1
.IC V(W_4_24_2) = 1 V(W_4_24_2_bar) = 0
.IC V(W_4_24_3) = 0 V(W_4_24_3_bar) = 1
.IC V(W_4_24_4) = 1 V(W_4_24_4_bar) = 0
.IC V(W_4_25_1) = 0 V(W_4_25_1_bar) = 1
.IC V(W_4_25_2) = 1 V(W_4_25_2_bar) = 0
.IC V(W_4_25_3) = 0 V(W_4_25_3_bar) = 1
.IC V(W_4_25_4) = 1 V(W_4_25_4_bar) = 0
.IC V(W_4_26_1) = 0 V(W_4_26_1_bar) = 1
.IC V(W_4_26_2) = 1 V(W_4_26_2_bar) = 0
.IC V(W_4_26_3) = 0 V(W_4_26_3_bar) = 1
.IC V(W_4_26_4) = 1 V(W_4_26_4_bar) = 0
.IC V(W_4_27_1) = 0 V(W_4_27_1_bar) = 1
.IC V(W_4_27_2) = 1 V(W_4_27_2_bar) = 0
.IC V(W_4_27_3) = 0 V(W_4_27_3_bar) = 1
.IC V(W_4_27_4) = 1 V(W_4_27_4_bar) = 0
.IC V(W_4_28_1) = 0 V(W_4_28_1_bar) = 1
.IC V(W_4_28_2) = 1 V(W_4_28_2_bar) = 0
.IC V(W_4_28_3) = 0 V(W_4_28_3_bar) = 1
.IC V(W_4_28_4) = 1 V(W_4_28_4_bar) = 0
.IC V(W_4_29_1) = 0 V(W_4_29_1_bar) = 1
.IC V(W_4_29_2) = 1 V(W_4_29_2_bar) = 0
.IC V(W_4_29_3) = 0 V(W_4_29_3_bar) = 1
.IC V(W_4_29_4) = 1 V(W_4_29_4_bar) = 0
.IC V(W_4_30_1) = 0 V(W_4_30_1_bar) = 1
.IC V(W_4_30_2) = 1 V(W_4_30_2_bar) = 0
.IC V(W_4_30_3) = 0 V(W_4_30_3_bar) = 1
.IC V(W_4_30_4) = 1 V(W_4_30_4_bar) = 0
.IC V(W_4_31_1) = 0 V(W_4_31_1_bar) = 1
.IC V(W_4_31_2) = 1 V(W_4_31_2_bar) = 0
.IC V(W_4_31_3) = 0 V(W_4_31_3_bar) = 1
.IC V(W_4_31_4) = 1 V(W_4_31_4_bar) = 0
.IC V(W_4_32_1) = 0 V(W_4_32_1_bar) = 1
.IC V(W_4_32_2) = 1 V(W_4_32_2_bar) = 0
.IC V(W_4_32_3) = 0 V(W_4_32_3_bar) = 1
.IC V(W_4_32_4) = 1 V(W_4_32_4_bar) = 0

.end
