.SUBCKT Control VSS VDD  clk rst_n out_valid
Xcounter_reg_0_ VSS VDD  clk N_8 n4 n13 n7 ASYNC_DFFHx1_ASAP7_75t_L
Xcounter_reg_2_ VSS VDD  clk N_10 n4 n8 n6 ASYNC_DFFHx1_ASAP7_75t_L
Xcounter_reg_1_ VSS VDD  clk N_9 n4 n12 n5 ASYNC_DFFHx1_ASAP7_75t_L
Xout_valid_reg VSS VDD   clk N_12 n4 n11 n3 ASYNC_DFFHx1_ASAP7_75t_L
XU12 VSS VDD  n7 n5 n9 NAND2xp33_ASAP7_75t_L
XU13 VSS VDD  n7 n5 n14 AND2x2_ASAP7_75t_L
XU14 VSS VDD  n6 n10 BUFx5_ASAP7_75t_L
XU15 VSS VDD  n10 n16 INVx3_ASAP7_75t_L
XU16 VSS VDD  rst_n n11 INVx6_ASAP7_75t_L
XU17 VSS VDD  rst_n n12 INVx6_ASAP7_75t_L
XU18 VSS VDD  rst_n n13 INVx6_ASAP7_75t_L
XU19 VSS VDD  rst_n n8 INVx6_ASAP7_75t_L
XU20 VSS VDD  n4 TIELOx1_ASAP7_75t_L
XU21 VSS VDD  n3 out_valid INVxp33_ASAP7_75t_L
XU22 VSS VDD  n10 n9 N_12 NOR2xp33_ASAP7_75t_L
XU23 VSS VDD  n7 n5 n15 NOR2xp33_ASAP7_75t_L
XU24 VSS VDD  n15 n16 n14 N_9 NOR3xp33_ASAP7_75t_L
XU25 VSS VDD  n10 n7 N_8 AND2x2_ASAP7_75t_L
XU26 VSS VDD  n7 n16 n5 N_10 NOR3xp33_ASAP7_75t_L
.ENDS


