.SUBCKT Control clk rst_n out_valid
Xcounter_reg_0_ N8 clk n4 n13 n7 ASYNC_DFFHx1_ASAP7_75t_R
Xcounter_reg_2_ N10 clk n4 n8 n6 ASYNC_DFFHx1_ASAP7_75t_R
Xcounter_reg_1_ N9 clk n4 n12 n5 ASYNC_DFFHx1_ASAP7_75t_R
Xout_valid_reg N12 clk n4 n11 n3 ASYNC_DFFHx1_ASAP7_75t_R
XU12 n6 n10 BUFx5_ASAP7_75t_R
XU13 n7 n5 n9 NAND2xp33_ASAP7_75t_R
XU14 n7 n5 n14 AND2x2_ASAP7_75t_R
XU15 n10 n16 INVx2_ASAP7_75t_R
XU16 rst_n n11 INVx8_ASAP7_75t_R
XU17 rst_n n12 INVx8_ASAP7_75t_R
XU18 rst_n n13 INVx8_ASAP7_75t_R
XU19 rst_n n8 INVx8_ASAP7_75t_R
XU20 n4 TIELOx1_ASAP7_75t_R
XU21 n3 out_valid INVxp33_ASAP7_75t_R
XU22 n10 n9 N12 NOR2xp33_ASAP7_75t_R
XU23 n7 n5 n15 NOR2xp33_ASAP7_75t_R
XU24 n15 n16 n14 N9 NOR3xp33_ASAP7_75t_R
XU25 n10 n7 N8 AND2x2_ASAP7_75t_R
XU26 n7 n16 n5 N10 NOR3xp33_ASAP7_75t_R
.ENDS


