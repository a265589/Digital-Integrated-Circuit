.SUBCKT Adder_tree VSS VDD  in[127] in[126] in[125] in[124] in[123] in[122] in[121] in[120] in[119] in[118] in[117] in[116] in[115] in[114] in[113] in[112] in[111] in[110] in[109] in[108] in[107] in[106] in[105] in[104] in[103] in[102] in[101] in[100] in[99] in[98] in[97] in[96] in[95] in[94] in[93] in[92] in[91] in[90] in[89] in[88] in[87] in[86] in[85] in[84] in[83] in[82] in[81] in[80] in[79] in[78] in[77] in[76] in[75] in[74] in[73] in[72] in[71] in[70] in[69] in[68] in[67] in[66] in[65] in[64] in[63] in[62] in[61] in[60] in[59] in[58] in[57] in[56] in[55] in[54] in[53] in[52] in[51] in[50] in[49] in[48] in[47] in[46] in[45] in[44] in[43] in[42] in[41] in[40] in[39] in[38] in[37] in[36] in[35] in[34] in[33] in[32] in[31] in[30] in[29] in[28] in[27] in[26] in[25] in[24] in[23] in[22] in[21] in[20] in[19] in[18] in[17] in[16] in[15] in[14] in[13] in[12] in[11] in[10] in[9] in[8] in[7] in[6] in[5] in[4] in[3] in[2] in[1] in[0] out[12] out[11] out[10] out[9] out[8] out[7] out[6] out[5] out[4] out[3] out[2] out[1] out[0]
XDP_OP_94J1_122_9915_U198 VSS VDD  in[4] in[28] in[36] DP_OP_94J1_122_9915_n299 DP_OP_94J1_122_9915_n300 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U197 VSS VDD  in[44] in[52] in[60] DP_OP_94J1_122_9915_n297 DP_OP_94J1_122_9915_n298 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U196 VSS VDD  in[68] in[76] in[84] DP_OP_94J1_122_9915_n295 DP_OP_94J1_122_9915_n296 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U195 VSS VDD  in[92] in[100] in[108] DP_OP_94J1_122_9915_n293 DP_OP_94J1_122_9915_n294 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U192 VSS VDD  in[88] in[80] in[72] DP_OP_94J1_122_9915_n287 DP_OP_94J1_122_9915_n288 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U190 VSS VDD  in[40] in[0] in[32] DP_OP_94J1_122_9915_n283 DP_OP_94J1_122_9915_n284 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U187 VSS VDD  DP_OP_94J1_122_9915_n286 DP_OP_94J1_122_9915_n278 DP_OP_94J1_122_9915_n284 DP_OP_94J1_122_9915_n279 DP_OP_94J1_122_9915_n280 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U186 VSS VDD  DP_OP_94J1_122_9915_n282 DP_OP_94J1_122_9915_n288 DP_OP_94J1_122_9915_n290 DP_OP_94J1_122_9915_n276 DP_OP_94J1_122_9915_n277 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U185 VSS VDD  DP_OP_94J1_122_9915_n292 DP_OP_94J1_122_9915_n294 DP_OP_94J1_122_9915_n296 DP_OP_94J1_122_9915_n274 DP_OP_94J1_122_9915_n275 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U183 VSS VDD  DP_OP_94J1_122_9915_n298 DP_OP_94J1_122_9915_n300 DP_OP_94J1_122_9915_n271 DP_OP_94J1_122_9915_n272 DP_OP_94J1_122_9915_n273 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U179 VSS VDD  in[45] in[53] in[61] DP_OP_94J1_122_9915_n265 DP_OP_94J1_122_9915_n266 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U178 VSS VDD  in[69] in[77] in[85] DP_OP_94J1_122_9915_n263 DP_OP_94J1_122_9915_n264 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U177 VSS VDD  in[93] in[101] in[109] DP_OP_94J1_122_9915_n261 DP_OP_94J1_122_9915_n262 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U174 VSS VDD  in[9] in[65] in[17] DP_OP_94J1_122_9915_n255 DP_OP_94J1_122_9915_n256 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U171 VSS VDD  in[57] in[41] in[49] DP_OP_94J1_122_9915_n249 DP_OP_94J1_122_9915_n250 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U169 VSS VDD  DP_OP_94J1_122_9915_n299 DP_OP_94J1_122_9915_n246 DP_OP_94J1_122_9915_n297 DP_OP_94J1_122_9915_n247 DP_OP_94J1_122_9915_n248 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U166 VSS VDD  DP_OP_94J1_122_9915_n285 DP_OP_94J1_122_9915_n281 DP_OP_94J1_122_9915_n287 DP_OP_94J1_122_9915_n241 DP_OP_94J1_122_9915_n242 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U165 VSS VDD  DP_OP_94J1_122_9915_n289 DP_OP_94J1_122_9915_n291 DP_OP_94J1_122_9915_n293 DP_OP_94J1_122_9915_n239 DP_OP_94J1_122_9915_n240 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U163 VSS VDD  DP_OP_94J1_122_9915_n258 n215 DP_OP_94J1_122_9915_n256 DP_OP_94J1_122_9915_n235 DP_OP_94J1_122_9915_n236 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U162 VSS VDD  DP_OP_94J1_122_9915_n266 DP_OP_94J1_122_9915_n254 DP_OP_94J1_122_9915_n264 DP_OP_94J1_122_9915_n233 DP_OP_94J1_122_9915_n234 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U156 VSS VDD  DP_OP_94J1_122_9915_n234 DP_OP_94J1_122_9915_n236 n100 DP_OP_94J1_122_9915_n224 DP_OP_94J1_122_9915_n225 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U148 VSS VDD  in[2] in[106] in[10] DP_OP_94J1_122_9915_n211 DP_OP_94J1_122_9915_n212 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U146 VSS VDD  in[86] in[26] in[34] DP_OP_94J1_122_9915_n207 DP_OP_94J1_122_9915_n208 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U143 VSS VDD  in[126] in[50] in[114] DP_OP_94J1_122_9915_n201 DP_OP_94J1_122_9915_n202 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U142 VSS VDD  in[58] in[90] in[66] DP_OP_94J1_122_9915_n199 DP_OP_94J1_122_9915_n200 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U141 VSS VDD  in[98] in[74] in[82] DP_OP_94J1_122_9915_n197 DP_OP_94J1_122_9915_n198 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U139 VSS VDD  DP_OP_94J1_122_9915_n267 DP_OP_94J1_122_9915_n194 DP_OP_94J1_122_9915_n265 DP_OP_94J1_122_9915_n195 DP_OP_94J1_122_9915_n196 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U137 VSS VDD  DP_OP_94J1_122_9915_n263 DP_OP_94J1_122_9915_n249 DP_OP_94J1_122_9915_n191 DP_OP_94J1_122_9915_n192 DP_OP_94J1_122_9915_n193 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U136 VSS VDD  DP_OP_94J1_122_9915_n251 DP_OP_94J1_122_9915_n257 DP_OP_94J1_122_9915_n261 DP_OP_94J1_122_9915_n189 DP_OP_94J1_122_9915_n190 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U135 VSS VDD  DP_OP_94J1_122_9915_n253 DP_OP_94J1_122_9915_n259 DP_OP_94J1_122_9915_n255 DP_OP_94J1_122_9915_n187 DP_OP_94J1_122_9915_n188 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U133 VSS VDD  DP_OP_94J1_122_9915_n247 DP_OP_94J1_122_9915_n241 n168 DP_OP_94J1_122_9915_n185 DP_OP_94J1_122_9915_n186 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U131 VSS VDD  DP_OP_94J1_122_9915_n210 DP_OP_94J1_122_9915_n202 n31 DP_OP_94J1_122_9915_n182 DP_OP_94J1_122_9915_n183 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U130 VSS VDD  DP_OP_94J1_122_9915_n214 DP_OP_94J1_122_9915_n204 DP_OP_94J1_122_9915_n216 DP_OP_94J1_122_9915_n179 DP_OP_94J1_122_9915_n180 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U125 VSS VDD  DP_OP_94J1_122_9915_n237 DP_OP_94J1_122_9915_n235 DP_OP_94J1_122_9915_n233 DP_OP_94J1_122_9915_n170 DP_OP_94J1_122_9915_n171 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U123 VSS VDD  DP_OP_94J1_122_9915_n228 DP_OP_94J1_122_9915_n231 DP_OP_94J1_122_9915_n167 DP_OP_94J1_122_9915_n168 DP_OP_94J1_122_9915_n169 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U113 VSS VDD  in[47] in[115] in[55] DP_OP_94J1_122_9915_n151 DP_OP_94J1_122_9915_n152 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U112 VSS VDD  in[63] in[3] in[71] DP_OP_94J1_122_9915_n149 DP_OP_94J1_122_9915_n150 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U111 VSS VDD  in[79] in[99] in[11] DP_OP_94J1_122_9915_n147 DP_OP_94J1_122_9915_n148 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U109 VSS VDD  in[95] in[27] in[103] DP_OP_94J1_122_9915_n143 DP_OP_94J1_122_9915_n144 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U106 VSS VDD  in[91] in[51] in[83] DP_OP_94J1_122_9915_n137 DP_OP_94J1_122_9915_n138 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U105 VSS VDD  in[75] in[59] in[67] DP_OP_94J1_122_9915_n135 DP_OP_94J1_122_9915_n136 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U101 VSS VDD  DP_OP_94J1_122_9915_n211 DP_OP_94J1_122_9915_n129 DP_OP_94J1_122_9915_n197 DP_OP_94J1_122_9915_n130 DP_OP_94J1_122_9915_n131 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U100 VSS VDD  DP_OP_94J1_122_9915_n209 n48 DP_OP_94J1_122_9915_n199 DP_OP_94J1_122_9915_n127 DP_OP_94J1_122_9915_n128 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U99 VSS VDD  DP_OP_94J1_122_9915_n207 DP_OP_94J1_122_9915_n203 DP_OP_94J1_122_9915_n201 DP_OP_94J1_122_9915_n125 DP_OP_94J1_122_9915_n126 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U93 VSS VDD  DP_OP_94J1_122_9915_n152 DP_OP_94J1_122_9915_n154 DP_OP_94J1_122_9915_n144 DP_OP_94J1_122_9915_n115 DP_OP_94J1_122_9915_n116 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U89 VSS VDD  n157 DP_OP_94J1_122_9915_n179 DP_OP_94J1_122_9915_n182 DP_OP_94J1_122_9915_n110 DP_OP_94J1_122_9915_n111 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U84 VSS VDD  DP_OP_94J1_122_9915_n124 n167 DP_OP_94J1_122_9915_n170 DP_OP_94J1_122_9915_n102 DP_OP_94J1_122_9915_n103 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U82 VSS VDD  DP_OP_94J1_122_9915_n172 DP_OP_94J1_122_9915_n114 n101 DP_OP_94J1_122_9915_n99 DP_OP_94J1_122_9915_n100 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U68 VSS VDD  DP_OP_94J1_122_9915_n147 DP_OP_94J1_122_9915_n143 DP_OP_94J1_122_9915_n135 DP_OP_94J1_122_9915_n78 DP_OP_94J1_122_9915_n79 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U66 VSS VDD  DP_OP_94J1_122_9915_n125 DP_OP_94J1_122_9915_n133 DP_OP_94J1_122_9915_n130 DP_OP_94J1_122_9915_n74 DP_OP_94J1_122_9915_n75 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U62 VSS VDD  DP_OP_94J1_122_9915_n81 DP_OP_94J1_122_9915_n117 DP_OP_94J1_122_9915_n79 DP_OP_94J1_122_9915_n67 DP_OP_94J1_122_9915_n68 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U61 VSS VDD  DP_OP_94J1_122_9915_n75 DP_OP_94J1_122_9915_n113 DP_OP_94J1_122_9915_n107 DP_OP_94J1_122_9915_n65 DP_OP_94J1_122_9915_n66 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U58 VSS VDD  DP_OP_94J1_122_9915_n71 DP_OP_94J1_122_9915_n68 n30 DP_OP_94J1_122_9915_n61 DP_OP_94J1_122_9915_n62 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U53 VSS VDD  DP_OP_94J1_122_9915_n76 DP_OP_94J1_122_9915_n83 DP_OP_94J1_122_9915_n80 DP_OP_94J1_122_9915_n51 DP_OP_94J1_122_9915_n52 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U50 VSS VDD  DP_OP_94J1_122_9915_n67 DP_OP_94J1_122_9915_n52 DP_OP_94J1_122_9915_n70 DP_OP_94J1_122_9915_n46 DP_OP_94J1_122_9915_n47 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U49 VSS VDD  DP_OP_94J1_122_9915_n50 DP_OP_94J1_122_9915_n65 DP_OP_94J1_122_9915_n63 DP_OP_94J1_122_9915_n44 DP_OP_94J1_122_9915_n45 FAx1_ASAP7_75t_L
XDP_OP_94J1_122_9915_U44 VSS VDD  DP_OP_94J1_122_9915_n46 DP_OP_94J1_122_9915_n49 n160 DP_OP_94J1_122_9915_n37 DP_OP_94J1_122_9915_n38 FAx1_ASAP7_75t_L
XU3 VSS VDD  DP_OP_94J1_122_9915_n37 n96 n197 XNOR2xp5_ASAP7_75t_L
XU4 VSS VDD  n129 n130 DP_OP_94J1_122_9915_n91 XOR2xp5_ASAP7_75t_L
XU5 VSS VDD  n147 DP_OP_94J1_122_9915_n227 n109 XNOR2xp5_ASAP7_75t_L
XU6 VSS VDD  n17 n153 n136 XOR2xp5_ASAP7_75t_L
XU7 VSS VDD  DP_OP_94J1_122_9915_n103 DP_OP_94J1_122_9915_n100 n130 XNOR2xp5_ASAP7_75t_L
XU8 VSS VDD  n174 n175 n108 XNOR2xp5_ASAP7_75t_L
XU9 VSS VDD  n91 n131 n90 XOR2xp5_ASAP7_75t_L
XU10 VSS VDD  n134 n65 n84 XNOR2xp5_ASAP7_75t_L
XU11 VSS VDD  n174 n175 n104 XOR2xp5_ASAP7_75t_L
XU12 VSS VDD  n193 n116 INVx1_ASAP7_75t_L
XU13 VSS VDD  n45 n91 INVx2_ASAP7_75t_L
XU14 VSS VDD  n57 n56 n44 XNOR2xp5_ASAP7_75t_L
XU15 VSS VDD  n154 n30 INVx2_ASAP7_75t_L
XU16 VSS VDD  DP_OP_94J1_122_9915_n123 n183 DP_OP_94J1_122_9915_n71 XOR2xp5_ASAP7_75t_L
XU17 VSS VDD  n176 n156 DP_OP_94J1_122_9915_n176 XNOR2xp5_ASAP7_75t_L
XU18 VSS VDD  n71 n70 DP_OP_94J1_122_9915_n227 XNOR2xp5_ASAP7_75t_L
XU19 VSS VDD  DP_OP_94J1_122_9915_n131 n16 n64 XNOR2xp5_ASAP7_75t_L
XU20 VSS VDD  n15 n37 n176 XNOR2xp5_ASAP7_75t_L
XU21 VSS VDD  n141 n140 n101 XNOR2xp5_ASAP7_75t_L
XU22 VSS VDD  in[7] in[15] DP_OP_94J1_122_9915_n129 XNOR2xp5_ASAP7_75t_L
XU23 VSS VDD  in[81] n88 n87 XNOR2xp5_ASAP7_75t_L
XU24 VSS VDD  in[117] in[1] n88 XOR2xp5_ASAP7_75t_L
XU25 VSS VDD  in[123] in[43] n139 XOR2xp5_ASAP7_75t_L
XU26 VSS VDD  DP_OP_94J1_122_9915_n198 n168 INVx1_ASAP7_75t_L
XU27 VSS VDD  n5 TIEHIx1_ASAP7_75t_L
XU28 VSS VDD  n5 out[9] INVx1_ASAP7_75t_L
XU29 VSS VDD  n5 out[10] INVx1_ASAP7_75t_L
XU30 VSS VDD  n5 out[11] INVx1_ASAP7_75t_L
XU31 VSS VDD  n5 out[12] INVx1_ASAP7_75t_L
XU32 VSS VDD  DP_OP_94J1_122_9915_n195 n6 DP_OP_94J1_122_9915_n124 XOR2xp5_ASAP7_75t_L
XU33 VSS VDD  n103 DP_OP_94J1_122_9915_n189 n6 XNOR2xp5_ASAP7_75t_L
XU34 VSS VDD  n63 n197 n32 n127 NAND3xp33_ASAP7_75t_L
XU35 VSS VDD  n51 n136 DP_OP_94J1_122_9915_n40 XNOR2xp5_ASAP7_75t_L
XU36 VSS VDD  DP_OP_94J1_122_9915_n102 n154 BUFx2_ASAP7_75t_L
XU37 VSS VDD  DP_OP_94J1_122_9915_n195 n103 DP_OP_94J1_122_9915_n189 n7 MAJIxp5_ASAP7_75t_L
XU38 VSS VDD  DP_OP_94J1_122_9915_n195 n103 DP_OP_94J1_122_9915_n189 DP_OP_94J1_122_9915_n123 MAJx2_ASAP7_75t_L
XU39 VSS VDD  n8 DP_OP_94J1_122_9915_n248 n100 XOR2x2_ASAP7_75t_L
XU40 VSS VDD  DP_OP_94J1_122_9915_n279 n47 n8 XOR2xp5_ASAP7_75t_L
XU41 VSS VDD  n55 n54 n32 AND2x2_ASAP7_75t_L
XU42 VSS VDD  in[14] in[6] DP_OP_94J1_122_9915_n132 NAND2xp5_ASAP7_75t_L
XU43 VSS VDD  n46 n123 n122 NAND2xp5_ASAP7_75t_L
XU44 VSS VDD  DP_OP_94J1_122_9915_n207 DP_OP_94J1_122_9915_n203 DP_OP_94J1_122_9915_n201 n9 MAJIxp5_ASAP7_75t_L
XU45 VSS VDD  n13 n29 n66 n10 MAJIxp5_ASAP7_75t_L
XU46 VSS VDD  n13 n29 n66 n11 MAJIxp5_ASAP7_75t_L
XU47 VSS VDD  DP_OP_94J1_122_9915_n200 DP_OP_94J1_122_9915_n206 DP_OP_94J1_122_9915_n212 n12 MAJIxp5_ASAP7_75t_L
XU48 VSS VDD  n129 n130 n13 XNOR2xp5_ASAP7_75t_L
XU49 VSS VDD  DP_OP_94J1_122_9915_n37 n96 n14 XOR2xp5_ASAP7_75t_L
XU50 VSS VDD  n34 DP_OP_94J1_122_9915_n283 DP_OP_94J1_122_9915_n295 n15 MAJIxp5_ASAP7_75t_L
XU51 VSS VDD  n34 DP_OP_94J1_122_9915_n283 DP_OP_94J1_122_9915_n295 DP_OP_94J1_122_9915_n244 MAJx2_ASAP7_75t_L
XU52 VSS VDD  DP_OP_94J1_122_9915_n200 DP_OP_94J1_122_9915_n206 DP_OP_94J1_122_9915_n212 n16 MAJx2_ASAP7_75t_L
XU53 VSS VDD  DP_OP_94J1_122_9915_n47 DP_OP_94J1_122_9915_n61 n17 XNOR2xp5_ASAP7_75t_L
XU54 VSS VDD  in[4] in[28] in[36] n18 MAJIxp5_ASAP7_75t_L
XU55 VSS VDD  n196 n98 n19 XOR2xp5_ASAP7_75t_L
XU56 VSS VDD  n196 n98 n59 XOR2xp5_ASAP7_75t_L
XU57 VSS VDD  DP_OP_94J1_122_9915_n226 DP_OP_94J1_122_9915_n176 n131 XOR2x2_ASAP7_75t_L
XU58 VSS VDD  n84 n193 n196 XNOR2x2_ASAP7_75t_L
XU59 VSS VDD  DP_OP_94J1_122_9915_n99 n118 BUFx4_ASAP7_75t_L
XU60 VSS VDD  DP_OP_94J1_122_9915_n168 n111 BUFx4_ASAP7_75t_L
XU61 VSS VDD  DP_OP_94J1_122_9915_n240 n25 BUFx4_ASAP7_75t_L
XU62 VSS VDD  in[30] in[38] in[22] n20 MAJIxp5_ASAP7_75t_L
XU63 VSS VDD  in[13] in[5] n21 XOR2xp5_ASAP7_75t_L
XU64 VSS VDD  n57 n56 n22 XOR2xp5_ASAP7_75t_L
XU65 VSS VDD  n60 n19 n23 XOR2xp5_ASAP7_75t_L
XU66 VSS VDD  DP_OP_94J1_122_9915_n245 n172 n24 XOR2xp5_ASAP7_75t_L
XU67 VSS VDD  in[81] n88 n26 XOR2xp5_ASAP7_75t_L
XU68 VSS VDD  n131 n45 n27 XNOR2xp5_ASAP7_75t_L
XU69 VSS VDD  n71 n70 n28 XOR2xp5_ASAP7_75t_L
XU70 VSS VDD  DP_OP_94J1_122_9915_n239 n159 BUFx4_ASAP7_75t_L
XU71 VSS VDD  n39 n73 INVx3_ASAP7_75t_L
XU72 VSS VDD  n78 DP_OP_94J1_122_9915_n161 n206 n29 MAJx2_ASAP7_75t_L
XU73 VSS VDD  n159 n31 INVx3_ASAP7_75t_L
XU74 VSS VDD  DP_OP_94J1_122_9915_n171 n45 BUFx4_ASAP7_75t_L
XU75 VSS VDD  in[13] in[5] n34 XNOR2xp5_ASAP7_75t_L
XU76 VSS VDD  n45 n131 n35 XOR2x2_ASAP7_75t_L
XU77 VSS VDD  DP_OP_94J1_122_9915_n183 n36 HB1xp67_ASAP7_75t_L
XU78 VSS VDD  n43 n170 HB1xp67_ASAP7_75t_L
XU79 VSS VDD  n170 n37 INVx1_ASAP7_75t_L
XU80 VSS VDD  n50 n163 n38 OR2x2_ASAP7_75t_L
XU81 VSS VDD  n37 n15 n102 NOR2xp33_ASAP7_75t_L
XU82 VSS VDD  n75 n39 BUFx6f_ASAP7_75t_L
XU83 VSS VDD  DP_OP_94J1_122_9915_n110 n76 n75 XNOR2x2_ASAP7_75t_L
XU84 VSS VDD  n78 n206 DP_OP_94J1_122_9915_n161 n40 MAJIxp5_ASAP7_75t_L
XU85 VSS VDD  DP_OP_94J1_122_9915_n245 n172 n41 XNOR2xp5_ASAP7_75t_L
XU86 VSS VDD  n60 n59 n42 XNOR2xp5_ASAP7_75t_L
XU87 VSS VDD  in[86] in[26] in[34] A0  n43 FAx1_ASAP7_75t_L
XU88 VSS VDD  n171 DP_OP_94J1_122_9915_n57 n42 n46 MAJIxp5_ASAP7_75t_L
XU89 VSS VDD  n121 n123 n63 NAND2xp33_ASAP7_75t_L
XU90 VSS VDD  DP_OP_94J1_122_9915_n244 DP_OP_94J1_122_9915_n208 n72 NOR2xp33_ASAP7_75t_L
XU91 VSS VDD  DP_OP_94J1_122_9915_n276 DP_OP_94J1_122_9915_n274 n69 NAND2xp33_ASAP7_75t_L
XU92 VSS VDD  in[13] in[5] DP_OP_94J1_122_9915_n194 NAND2xp5_ASAP7_75t_L
XU93 VSS VDD  n69 n71 n68 NAND2xp33_ASAP7_75t_L
XU94 VSS VDD  in[7] in[15] n213 NAND2xp33_ASAP7_75t_L
XU95 VSS VDD  DP_OP_94J1_122_9915_n77 DP_OP_94J1_122_9915_n120 n183 XNOR2xp5_ASAP7_75t_L
XU96 VSS VDD  in[21] n62 n47 XOR2xp5_ASAP7_75t_L
XU97 VSS VDD  in[122] in[102] in[94] n48 MAJIxp5_ASAP7_75t_L
XU98 VSS VDD  DP_OP_94J1_122_9915_n276 DP_OP_94J1_122_9915_n274 n49 OR2x2_ASAP7_75t_L
XU99 VSS VDD  DP_OP_94J1_122_9915_n56 DP_OP_94J1_122_9915_n45 n136 n50 MAJIxp5_ASAP7_75t_L
XU100 VSS VDD  in[127] n139 n103 XOR2xp5_ASAP7_75t_L
XU101 VSS VDD  n14 n38 n126 AND2x2_ASAP7_75t_L
XU102 VSS VDD  n111 n155 INVx2_ASAP7_75t_L
XU103 VSS VDD  n118 n134 INVx2_ASAP7_75t_L
XU104 VSS VDD  n162 n161 INVx2_ASAP7_75t_L
XU105 VSS VDD  n117 n65 INVxp67_ASAP7_75t_L
XU106 VSS VDD  n102 n135 n57 NOR2xp67_ASAP7_75t_L
XU107 VSS VDD  n72 n115 n135 NOR2xp33_ASAP7_75t_L
XU108 VSS VDD  DP_OP_94J1_122_9915_n196 n156 INVxp67_ASAP7_75t_L
XU109 VSS VDD  n25 n173 INVx2_ASAP7_75t_L
XU110 VSS VDD  DP_OP_94J1_122_9915_n200 n177 DP_OP_94J1_122_9915_n178 XOR2xp5_ASAP7_75t_L
XU111 VSS VDD  in[38] in[30] n133 XOR2xp5_ASAP7_75t_L
XU112 VSS VDD  n210 DP_OP_94J1_122_9915_n40 n123 OR2x2_ASAP7_75t_L
XU113 VSS VDD  n116 DP_OP_94J1_122_9915_n66 n118 n153 MAJx2_ASAP7_75t_L
XU114 VSS VDD  DP_OP_94J1_122_9915_n56 n52 n51 XNOR2xp5_ASAP7_75t_L
XU115 VSS VDD  n114 n52 INVxp67_ASAP7_75t_L
XU116 VSS VDD  DP_OP_94J1_122_9915_n62 n53 n73 DP_OP_94J1_122_9915_n56 MAJIxp5_ASAP7_75t_L
XU117 VSS VDD  n125 n127 n158 out[7] NAND3xp33_ASAP7_75t_L
XU118 VSS VDD  n53 n39 n74 XNOR2xp5_ASAP7_75t_L
XU119 VSS VDD  DP_OP_94J1_122_9915_n162 n44 n216 n53 MAJIxp5_ASAP7_75t_L
XU120 VSS VDD  n163 n50 n54 NAND2xp5_ASAP7_75t_L
XU121 VSS VDD  n210 DP_OP_94J1_122_9915_n40 n55 NAND2xp5_ASAP7_75t_L
XU122 VSS VDD  DP_OP_94J1_122_9915_n116 DP_OP_94J1_122_9915_n126 n57 DP_OP_94J1_122_9915_n105 MAJIxp5_ASAP7_75t_L
XU123 VSS VDD  DP_OP_94J1_122_9915_n126 DP_OP_94J1_122_9915_n116 n56 XOR2xp5_ASAP7_75t_L
XU124 VSS VDD  DP_OP_94J1_122_9915_n193 DP_OP_94J1_122_9915_n188 DP_OP_94J1_122_9915_n190 DP_OP_94J1_122_9915_n172 MAJIxp5_ASAP7_75t_L
XU125 VSS VDD  DP_OP_94J1_122_9915_n193 n58 DP_OP_94J1_122_9915_n173 XOR2xp5_ASAP7_75t_L
XU126 VSS VDD  DP_OP_94J1_122_9915_n188 DP_OP_94J1_122_9915_n190 n58 XNOR2xp5_ASAP7_75t_L
XU127 VSS VDD  n13 n29 n66 n171 MAJIxp5_ASAP7_75t_L
XU128 VSS VDD  n195 n61 n66 XNOR2xp5_ASAP7_75t_L
XU129 VSS VDD  n10 DP_OP_94J1_122_9915_n57 n42 n121 MAJIxp5_ASAP7_75t_L
XU130 VSS VDD  n194 n195 n108 n60 MAJIxp5_ASAP7_75t_L
XU131 VSS VDD  n104 n194 n61 XOR2xp5_ASAP7_75t_L
XU132 VSS VDD  in[21] in[37] in[29] DP_OP_94J1_122_9915_n267 MAJIxp5_ASAP7_75t_L
XU133 VSS VDD  in[37] in[29] n62 XOR2xp5_ASAP7_75t_L
XU134 VSS VDD  DP_OP_94J1_122_9915_n128 DP_OP_94J1_122_9915_n131 n12 DP_OP_94J1_122_9915_n107 MAJIxp5_ASAP7_75t_L
XU135 VSS VDD  DP_OP_94J1_122_9915_n128 n64 DP_OP_94J1_122_9915_n108 XNOR2xp5_ASAP7_75t_L
XU136 VSS VDD  n66 DP_OP_94J1_122_9915_n91 n208 XNOR2xp5_ASAP7_75t_L
XU137 VSS VDD  n67 n27 n78 XNOR2xp5_ASAP7_75t_L
XU138 VSS VDD  n35 n67 n205 XNOR2xp5_ASAP7_75t_L
XU139 VSS VDD  DP_OP_94J1_122_9915_n169 DP_OP_94J1_122_9915_n221 n67 XNOR2xp5_ASAP7_75t_L
XU140 VSS VDD  n49 n68 DP_OP_94J1_122_9915_n226 NAND2xp5_ASAP7_75t_L
XU141 VSS VDD  DP_OP_94J1_122_9915_n274 DP_OP_94J1_122_9915_n276 n70 XNOR2xp5_ASAP7_75t_L
XU142 VSS VDD  n81 n26 n71 XOR2xp5_ASAP7_75t_L
XU143 VSS VDD  n74 DP_OP_94J1_122_9915_n62 DP_OP_94J1_122_9915_n57 XNOR2xp5_ASAP7_75t_L
XU144 VSS VDD  DP_OP_94J1_122_9915_n73 DP_OP_94J1_122_9915_n105 n76 XNOR2xp5_ASAP7_75t_L
XU145 VSS VDD  n45 DP_OP_94J1_122_9915_n226 DP_OP_94J1_122_9915_n176 DP_OP_94J1_122_9915_n162 MAJx2_ASAP7_75t_L
XU146 VSS VDD  n77 DP_OP_94J1_122_9915_n225 n204 n206 MAJIxp5_ASAP7_75t_L
XU147 VSS VDD  n147 n28 n77 XNOR2xp5_ASAP7_75t_L
XU148 VSS VDD  n24 n107 n147 XNOR2xp5_ASAP7_75t_L
XU149 VSS VDD  n107 n41 DP_OP_94J1_122_9915_n227 DP_OP_94J1_122_9915_n221 MAJIxp5_ASAP7_75t_L
XU150 VSS VDD  n80 n79 DP_OP_94J1_122_9915_n50 XNOR2xp5_ASAP7_75t_L
XU151 VSS VDD  n166 DP_OP_94J1_122_9915_n74 n79 XOR2xp5_ASAP7_75t_L
XU152 VSS VDD  n166 n80 DP_OP_94J1_122_9915_n74 DP_OP_94J1_122_9915_n49 MAJIxp5_ASAP7_75t_L
XU153 VSS VDD  DP_OP_94J1_122_9915_n115 DP_OP_94J1_122_9915_n84 DP_OP_94J1_122_9915_n127 n80 MAJIxp5_ASAP7_75t_L
XU154 VSS VDD  DP_OP_94J1_122_9915_n250 DP_OP_94J1_122_9915_n262 n81 XNOR2xp5_ASAP7_75t_L
XU155 VSS VDD  n20 DP_OP_94J1_122_9915_n213 DP_OP_94J1_122_9915_n132 DP_OP_94J1_122_9915_n133 MAJIxp5_ASAP7_75t_L
XU156 VSS VDD  n83 n82 DP_OP_94J1_122_9915_n134 XNOR2xp5_ASAP7_75t_L
XU157 VSS VDD  DP_OP_94J1_122_9915_n132 DP_OP_94J1_122_9915_n213 n82 XNOR2xp5_ASAP7_75t_L
XU158 VSS VDD  in[30] in[38] in[22] n83 MAJx2_ASAP7_75t_L
XU159 VSS VDD  n120 n119 n163 XNOR2xp5_ASAP7_75t_L
XU160 VSS VDD  n179 n85 n178 NAND2xp33_ASAP7_75t_L
XU161 VSS VDD  n126 n85 n125 NAND2xp5_ASAP7_75t_L
XU162 VSS VDD  n122 n32 n85 NAND2xp5_ASAP7_75t_L
XU163 VSS VDD  n86 n21 DP_OP_94J1_122_9915_n245 XNOR2xp5_ASAP7_75t_L
XU164 VSS VDD  DP_OP_94J1_122_9915_n283 DP_OP_94J1_122_9915_n295 n86 XNOR2xp5_ASAP7_75t_L
XU165 VSS VDD  DP_OP_94J1_122_9915_n262 n87 DP_OP_94J1_122_9915_n250 DP_OP_94J1_122_9915_n237 MAJIxp5_ASAP7_75t_L
XU166 VSS VDD  DP_OP_94J1_122_9915_n162 n89 n194 XNOR2xp5_ASAP7_75t_L
XU167 VSS VDD  n216 n22 n89 XNOR2xp5_ASAP7_75t_L
XU168 VSS VDD  DP_OP_94J1_122_9915_n169 n90 DP_OP_94J1_122_9915_n221 n195 MAJx2_ASAP7_75t_L
XU169 VSS VDD  n212 n92 out[6] XOR2xp5_ASAP7_75t_L
XU170 VSS VDD  DP_OP_94J1_122_9915_n40 n210 n121 n92 MAJIxp5_ASAP7_75t_L
XU171 VSS VDD  n9 DP_OP_94J1_122_9915_n133 DP_OP_94J1_122_9915_n130 A1  n93 FAx1_ASAP7_75t_L
XU172 VSS VDD  in[45] in[53] in[61] n94 MAJIxp5_ASAP7_75t_L
XU173 VSS VDD  n97 DP_OP_94J1_122_9915_n37 n180 NAND2xp33_ASAP7_75t_L
XU174 VSS VDD  in[78] in[18] n192 XOR2xp5_ASAP7_75t_L
XU175 VSS VDD  in[102] in[122] n201 XOR2xp5_ASAP7_75t_L
XU176 VSS VDD  in[16] in[8] n198 XOR2xp5_ASAP7_75t_L
XU177 VSS VDD  DP_OP_94J1_122_9915_n37 n97 n164 OR2x2_ASAP7_75t_L
XU178 VSS VDD  n129 DP_OP_94J1_122_9915_n103 DP_OP_94J1_122_9915_n100 n95 MAJIxp5_ASAP7_75t_L
XU179 VSS VDD  n120 DP_OP_94J1_122_9915_n44 DP_OP_94J1_122_9915_n38 n96 MAJIxp5_ASAP7_75t_L
XU180 VSS VDD  n111 DP_OP_94J1_122_9915_n108 n174 XOR2x2_ASAP7_75t_L
XU181 VSS VDD  n155 DP_OP_94J1_122_9915_n108 n151 n193 MAJx3_ASAP7_75t_L
XU182 VSS VDD  n120 DP_OP_94J1_122_9915_n44 DP_OP_94J1_122_9915_n38 n97 MAJx2_ASAP7_75t_L
XU183 VSS VDD  n129 DP_OP_94J1_122_9915_n103 DP_OP_94J1_122_9915_n100 n98 MAJx2_ASAP7_75t_L
XU184 VSS VDD  DP_OP_94J1_122_9915_n187 n105 BUFx4_ASAP7_75t_L
XU185 VSS VDD  DP_OP_94J1_122_9915_n272 n148 BUFx4_ASAP7_75t_L
XU186 VSS VDD  in[35] in[119] in[111] n99 MAJIxp5_ASAP7_75t_L
XU187 VSS VDD  DP_OP_94J1_122_9915_n136 DP_OP_94J1_122_9915_n150 n140 XNOR2x2_ASAP7_75t_L
XU188 VSS VDD  in[63] in[3] in[71] n110 MAJx2_ASAP7_75t_L
XU189 VSS VDD  DP_OP_94J1_122_9915_n209 n48 DP_OP_94J1_122_9915_n199 n113 MAJx2_ASAP7_75t_L
XU190 VSS VDD  n105 n141 INVx3_ASAP7_75t_L
XU191 VSS VDD  DP_OP_94J1_122_9915_n280 n106 HB1xp67_ASAP7_75t_L
XU192 VSS VDD  n148 n107 INVx3_ASAP7_75t_L
XU193 VSS VDD  n18 DP_OP_94J1_122_9915_n246 DP_OP_94J1_122_9915_n297 A2  n112 FAx1_ASAP7_75t_L
XU194 VSS VDD  DP_OP_94J1_122_9915_n50 DP_OP_94J1_122_9915_n65 DP_OP_94J1_122_9915_n63 A3  n114 FAx1_ASAP7_75t_L
XU195 VSS VDD  DP_OP_94J1_122_9915_n267 DP_OP_94J1_122_9915_n194 n94 A4  n115 FAx1_ASAP7_75t_L
XU196 VSS VDD  n93 DP_OP_94J1_122_9915_n113 DP_OP_94J1_122_9915_n107 A5  n117 FAx1_ASAP7_75t_L
XU197 VSS VDD  n112 n47 DP_OP_94J1_122_9915_n279 DP_OP_94J1_122_9915_n231 MAJIxp5_ASAP7_75t_L
XU198 VSS VDD  DP_OP_94J1_122_9915_n44 DP_OP_94J1_122_9915_n38 n119 XOR2xp5_ASAP7_75t_L
XU199 VSS VDD  n153 DP_OP_94J1_122_9915_n47 DP_OP_94J1_122_9915_n61 n120 MAJIxp5_ASAP7_75t_L
XU200 VSS VDD  in[64] in[48] in[56] DP_OP_94J1_122_9915_n285 MAJIxp5_ASAP7_75t_L
XU201 VSS VDD  in[64] n124 DP_OP_94J1_122_9915_n286 XNOR2xp5_ASAP7_75t_L
XU202 VSS VDD  in[48] in[56] n124 XOR2xp5_ASAP7_75t_L
XU203 VSS VDD  in[46] in[62] in[54] DP_OP_94J1_122_9915_n213 MAJIxp5_ASAP7_75t_L
XU204 VSS VDD  in[46] n128 DP_OP_94J1_122_9915_n214 XNOR2xp5_ASAP7_75t_L
XU205 VSS VDD  in[62] in[54] n128 XOR2xp5_ASAP7_75t_L
XU206 VSS VDD  DP_OP_94J1_122_9915_n224 DP_OP_94J1_122_9915_n173 n186 n129 MAJIxp5_ASAP7_75t_L
XU207 VSS VDD  DP_OP_94J1_122_9915_n273 DP_OP_94J1_122_9915_n275 DP_OP_94J1_122_9915_n277 n204 MAJIxp5_ASAP7_75t_L
XU208 VSS VDD  in[113] in[25] in[97] DP_OP_94J1_122_9915_n253 MAJIxp5_ASAP7_75t_L
XU209 VSS VDD  in[113] n132 DP_OP_94J1_122_9915_n254 XNOR2xp5_ASAP7_75t_L
XU210 VSS VDD  in[25] in[97] n132 XOR2xp5_ASAP7_75t_L
XU211 VSS VDD  in[22] n133 DP_OP_94J1_122_9915_n216 XNOR2xp5_ASAP7_75t_L
XU212 VSS VDD  n99 DP_OP_94J1_122_9915_n139 DP_OP_94J1_122_9915_n145 DP_OP_94J1_122_9915_n76 MAJIxp5_ASAP7_75t_L
XU213 VSS VDD  n138 n137 DP_OP_94J1_122_9915_n77 XNOR2xp5_ASAP7_75t_L
XU214 VSS VDD  DP_OP_94J1_122_9915_n139 DP_OP_94J1_122_9915_n145 n137 XNOR2xp5_ASAP7_75t_L
XU215 VSS VDD  in[35] in[119] in[111] n138 MAJx2_ASAP7_75t_L
XU216 VSS VDD  in[127] in[123] in[43] DP_OP_94J1_122_9915_n139 MAJIxp5_ASAP7_75t_L
XU217 VSS VDD  n141 DP_OP_94J1_122_9915_n136 DP_OP_94J1_122_9915_n150 DP_OP_94J1_122_9915_n120 MAJIxp5_ASAP7_75t_L
XU218 VSS VDD  DP_OP_94J1_122_9915_n149 DP_OP_94J1_122_9915_n137 DP_OP_94J1_122_9915_n151 DP_OP_94J1_122_9915_n80 MAJIxp5_ASAP7_75t_L
XU219 VSS VDD  n110 n142 DP_OP_94J1_122_9915_n81 XNOR2xp5_ASAP7_75t_L
XU220 VSS VDD  DP_OP_94J1_122_9915_n137 DP_OP_94J1_122_9915_n151 n142 XNOR2xp5_ASAP7_75t_L
XU221 VSS VDD  in[23] in[39] in[31] DP_OP_94J1_122_9915_n153 MAJIxp5_ASAP7_75t_L
XU222 VSS VDD  in[23] n143 DP_OP_94J1_122_9915_n154 XNOR2xp5_ASAP7_75t_L
XU223 VSS VDD  in[39] in[31] n143 XOR2xp5_ASAP7_75t_L
XU224 VSS VDD  n144 DP_OP_94J1_122_9915_n115 DP_OP_94J1_122_9915_n73 XNOR2xp5_ASAP7_75t_L
XU225 VSS VDD  n113 DP_OP_94J1_122_9915_n84 n144 XNOR2xp5_ASAP7_75t_L
XU226 VSS VDD  in[19] in[87] in[107] DP_OP_94J1_122_9915_n145 MAJIxp5_ASAP7_75t_L
XU227 VSS VDD  in[19] n145 DP_OP_94J1_122_9915_n146 XNOR2xp5_ASAP7_75t_L
XU228 VSS VDD  in[87] in[107] n145 XOR2xp5_ASAP7_75t_L
XU229 VSS VDD  in[125] in[121] in[89] DP_OP_94J1_122_9915_n257 MAJIxp5_ASAP7_75t_L
XU230 VSS VDD  in[125] n146 DP_OP_94J1_122_9915_n258 XNOR2xp5_ASAP7_75t_L
XU231 VSS VDD  in[121] in[89] n146 XOR2xp5_ASAP7_75t_L
XU232 VSS VDD  n164 n178 out[8] NAND2xp33_ASAP7_75t_L
XU233 VSS VDD  n194 n108 n195 n149 MAJIxp5_ASAP7_75t_L
XU234 VSS VDD  in[58] in[90] in[66] A6  n150 FAx1_ASAP7_75t_L
XU235 VSS VDD  DP_OP_94J1_122_9915_n111 n151 BUFx4_ASAP7_75t_L
XU236 VSS VDD  n150 n177 n152 XNOR2xp5_ASAP7_75t_L
XU237 VSS VDD  n163 n50 n212 XNOR2xp5_ASAP7_75t_L
XU238 VSS VDD  DP_OP_94J1_122_9915_n185 DP_OP_94J1_122_9915_n109 BUFx4_ASAP7_75t_L
XU239 VSS VDD  n151 n175 INVx3_ASAP7_75t_L
XU240 VSS VDD  DP_OP_94J1_122_9915_n109 n157 INVx3_ASAP7_75t_L
XU241 VSS VDD  DP_OP_94J1_122_9915_n186 n162 BUFx4_ASAP7_75t_L
XU242 VSS VDD  n106 DP_OP_94J1_122_9915_n271 INVx1_ASAP7_75t_L
XU243 VSS VDD  n38 n180 n179 AND2x2_ASAP7_75t_L
XU244 VSS VDD  n14 n38 n158 OR2x2_ASAP7_75t_L
XU245 VSS VDD  DP_OP_94J1_122_9915_n51 DP_OP_94J1_122_9915_n36 BUFx4_ASAP7_75t_L
XU246 VSS VDD  DP_OP_94J1_122_9915_n36 n160 INVx3_ASAP7_75t_L
XU247 VSS VDD  DP_OP_94J1_122_9915_n138 n199 BUFx4_ASAP7_75t_L
XU248 VSS VDD  n36 DP_OP_94J1_122_9915_n167 INVx1_ASAP7_75t_L
XU249 VSS VDD  DP_OP_94J1_122_9915_n78 DP_OP_94J1_122_9915_n48 BUFx4_ASAP7_75t_L
XU250 VSS VDD  DP_OP_94J1_122_9915_n153 n213 DP_OP_94J1_122_9915_n83 NOR2x1_ASAP7_75t_L
XU251 VSS VDD  DP_OP_94J1_122_9915_n120 DP_OP_94J1_122_9915_n77 n165 OR2x2_ASAP7_75t_L
XU252 VSS VDD  DP_OP_94J1_122_9915_n48 n166 INVx3_ASAP7_75t_L
XU253 VSS VDD  DP_OP_94J1_122_9915_n146 n191 n167 XNOR2xp5_ASAP7_75t_L
XU254 VSS VDD  n199 n169 INVx3_ASAP7_75t_L
XU255 VSS VDD  n25 DP_OP_94J1_122_9915_n242 DP_OP_94J1_122_9915_n245 DP_OP_94J1_122_9915_n228 MAJIxp5_ASAP7_75t_L
XU256 VSS VDD  DP_OP_94J1_122_9915_n242 n173 n172 XNOR2xp5_ASAP7_75t_L
XU257 VSS VDD  n210 DP_OP_94J1_122_9915_n40 n211 XNOR2xp5_ASAP7_75t_L
XU258 VSS VDD  DP_OP_94J1_122_9915_n206 DP_OP_94J1_122_9915_n212 n177 XNOR2xp5_ASAP7_75t_L
XU259 VSS VDD  n181 n165 DP_OP_94J1_122_9915_n70 NAND2xp5_ASAP7_75t_L
XU260 VSS VDD  n7 n182 n181 NAND2xp33_ASAP7_75t_L
XU261 VSS VDD  DP_OP_94J1_122_9915_n77 DP_OP_94J1_122_9915_n120 n182 NAND2xp5_ASAP7_75t_L
XU262 VSS VDD  in[111] n184 DP_OP_94J1_122_9915_n142 XNOR2xp5_ASAP7_75t_L
XU263 VSS VDD  in[119] in[35] n184 XOR2xp5_ASAP7_75t_L
XU264 VSS VDD  DP_OP_94J1_122_9915_n224 n185 DP_OP_94J1_122_9915_n161 XNOR2xp5_ASAP7_75t_L
XU265 VSS VDD  n186 DP_OP_94J1_122_9915_n173 n185 XOR2xp5_ASAP7_75t_L
XU266 VSS VDD  n187 n162 n186 XNOR2xp5_ASAP7_75t_L
XU267 VSS VDD  DP_OP_94J1_122_9915_n180 n152 n187 XOR2xp5_ASAP7_75t_L
XU268 VSS VDD  in[112] in[96] in[104] DP_OP_94J1_122_9915_n289 MAJIxp5_ASAP7_75t_L
XU269 VSS VDD  in[112] n188 DP_OP_94J1_122_9915_n290 XNOR2xp5_ASAP7_75t_L
XU270 VSS VDD  in[96] in[104] n188 XOR2xp5_ASAP7_75t_L
XU271 VSS VDD  DP_OP_94J1_122_9915_n110 DP_OP_94J1_122_9915_n73 DP_OP_94J1_122_9915_n105 DP_OP_94J1_122_9915_n63 MAJIxp5_ASAP7_75t_L
XU272 VSS VDD  in[110] in[118] in[42] DP_OP_94J1_122_9915_n203 MAJIxp5_ASAP7_75t_L
XU273 VSS VDD  in[110] n189 DP_OP_94J1_122_9915_n204 XNOR2xp5_ASAP7_75t_L
XU274 VSS VDD  in[118] in[42] n189 XOR2xp5_ASAP7_75t_L
XU275 VSS VDD  in[116] in[120] in[124] DP_OP_94J1_122_9915_n291 MAJIxp5_ASAP7_75t_L
XU276 VSS VDD  in[116] n190 DP_OP_94J1_122_9915_n292 XNOR2xp5_ASAP7_75t_L
XU277 VSS VDD  in[120] in[124] n190 XOR2xp5_ASAP7_75t_L
XU278 VSS VDD  DP_OP_94J1_122_9915_n146 DP_OP_94J1_122_9915_n142 DP_OP_94J1_122_9915_n148 DP_OP_94J1_122_9915_n117 MAJIxp5_ASAP7_75t_L
XU279 VSS VDD  DP_OP_94J1_122_9915_n142 DP_OP_94J1_122_9915_n148 n191 XNOR2xp5_ASAP7_75t_L
XU280 VSS VDD  in[70] in[78] in[18] DP_OP_94J1_122_9915_n209 MAJIxp5_ASAP7_75t_L
XU281 VSS VDD  in[70] n192 DP_OP_94J1_122_9915_n210 XNOR2xp5_ASAP7_75t_L
XU282 VSS VDD  in[20] in[12] DP_OP_94J1_122_9915_n246 NAND2xp5_ASAP7_75t_L
XU283 VSS VDD  n161 DP_OP_94J1_122_9915_n178 DP_OP_94J1_122_9915_n180 n216 MAJIxp5_ASAP7_75t_L
XU284 VSS VDD  n196 n95 n149 n210 MAJIxp5_ASAP7_75t_L
XU285 VSS VDD  in[105] in[73] in[33] DP_OP_94J1_122_9915_n251 MAJIxp5_ASAP7_75t_L
XU286 VSS VDD  in[24] in[16] in[8] DP_OP_94J1_122_9915_n281 MAJIxp5_ASAP7_75t_L
XU287 VSS VDD  in[24] n198 DP_OP_94J1_122_9915_n282 XNOR2xp5_ASAP7_75t_L
XU288 VSS VDD  n169 DP_OP_94J1_122_9915_n192 DP_OP_94J1_122_9915_n134 DP_OP_94J1_122_9915_n113 MAJIxp5_ASAP7_75t_L
XU289 VSS VDD  DP_OP_94J1_122_9915_n192 n169 n200 XNOR2xp5_ASAP7_75t_L
XU290 VSS VDD  DP_OP_94J1_122_9915_n134 n200 DP_OP_94J1_122_9915_n114 XOR2xp5_ASAP7_75t_L
XU291 VSS VDD  in[94] n201 DP_OP_94J1_122_9915_n206 XNOR2xp5_ASAP7_75t_L
XU292 VSS VDD  in[117] in[1] in[81] DP_OP_94J1_122_9915_n259 MAJIxp5_ASAP7_75t_L
XU293 VSS VDD  in[14] in[6] A7  DP_OP_94J1_122_9915_n191 HAxp5_ASAP7_75t_L
XU294 VSS VDD  in[20] in[12] A8  DP_OP_94J1_122_9915_n278 HAxp5_ASAP7_75t_L
XU295 VSS VDD  DP_OP_94J1_122_9915_n277 DP_OP_94J1_122_9915_n275 A9  n202 HAxp5_ASAP7_75t_L
XU296 VSS VDD  DP_OP_94J1_122_9915_n273 n202 A10  out[0] HAxp5_ASAP7_75t_L
XU297 VSS VDD  DP_OP_94J1_122_9915_n225 n109 A11  n203 HAxp5_ASAP7_75t_L
XU298 VSS VDD  n204 n203 A12  out[1] HAxp5_ASAP7_75t_L
XU299 VSS VDD  DP_OP_94J1_122_9915_n161 n205 n207 XOR2xp5_ASAP7_75t_L
XU300 VSS VDD  n207 n206 A13  out[2] HAxp5_ASAP7_75t_L
XU301 VSS VDD  n208 n40 A14  out[3] HAxp5_ASAP7_75t_L
XU302 VSS VDD  DP_OP_94J1_122_9915_n57 n23 A15  n209 HAxp5_ASAP7_75t_L
XU303 VSS VDD  n209 n11 A16  out[4] HAxp5_ASAP7_75t_L
XU304 VSS VDD  n211 n46 A17  out[5] HAxp5_ASAP7_75t_L
XU305 VSS VDD  DP_OP_94J1_122_9915_n153 n213 DP_OP_94J1_122_9915_n84 XOR2xp5_ASAP7_75t_L
XU306 VSS VDD  in[73] in[33] n214 XOR2xp5_ASAP7_75t_L
XU307 VSS VDD  in[105] n214 n215 XNOR2xp5_ASAP7_75t_L
.ENDS


