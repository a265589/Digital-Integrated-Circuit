.SUBCKT Adder_tree in[127] in[126] in[125] in[124] in[123] in[122] in[121] in[120] in[119] in[118] in[117] in[116] in[115] in[114] in[113] in[112] in[111] in[110] in[109] in[108] in[107] in[106] in[105] in[104] in[103] in[102] in[101] in[100] in[99] in[98] in[97] in[96] in[95] in[94] in[93] in[92] in[91] in[90] in[89] in[88] in[87] in[86] in[85] in[84] in[83] in[82] in[81] in[80] in[79] in[78] in[77] in[76] in[75] in[74] in[73] in[72] in[71] in[70] in[69] in[68] in[67] in[66] in[65] in[64] in[63] in[62] in[61] in[60] in[59] in[58] in[57] in[56] in[55] in[54] in[53] in[52] in[51] in[50] in[49] in[48] in[47] in[46] in[45] in[44] in[43] in[42] in[41] in[40] in[39] in[38] in[37] in[36] in[35] in[34] in[33] in[32] in[31] in[30] in[29] in[28] in[27] in[26] in[25] in[24] in[23] in[22] in[21] in[20] in[19] in[18] in[17] in[16] in[15] in[14] in[13] in[12] in[11] in[10] in[9] in[8] in[7] in[6] in[5] in[4] in[3] in[2] in[1] in[0] out[12] out[11] out[10] out[9] out[8] out[7] out[6] out[5] out[4] out[3] out[2] out[1] out[0]
XDP_OP_94J1_122_9915_U198 in[4] in[28] in[36] DP_OP_94J1_122_9915_n299 DP_OP_94J1_122_9915_n300 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U197 in[44] in[52] in[60] DP_OP_94J1_122_9915_n297 DP_OP_94J1_122_9915_n298 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U196 in[68] in[76] in[84] DP_OP_94J1_122_9915_n295 DP_OP_94J1_122_9915_n296 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U195 in[92] in[100] in[108] DP_OP_94J1_122_9915_n293 DP_OP_94J1_122_9915_n294 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U192 in[88] in[80] in[72] DP_OP_94J1_122_9915_n287 DP_OP_94J1_122_9915_n288 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U190 in[40] in[0] in[32] DP_OP_94J1_122_9915_n283 DP_OP_94J1_122_9915_n284 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U187 DP_OP_94J1_122_9915_n286 DP_OP_94J1_122_9915_n278 DP_OP_94J1_122_9915_n284 DP_OP_94J1_122_9915_n279 DP_OP_94J1_122_9915_n280 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U186 DP_OP_94J1_122_9915_n282 DP_OP_94J1_122_9915_n288 DP_OP_94J1_122_9915_n290 DP_OP_94J1_122_9915_n276 DP_OP_94J1_122_9915_n277 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U185 DP_OP_94J1_122_9915_n292 DP_OP_94J1_122_9915_n294 DP_OP_94J1_122_9915_n296 DP_OP_94J1_122_9915_n274 DP_OP_94J1_122_9915_n275 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U183 DP_OP_94J1_122_9915_n298 DP_OP_94J1_122_9915_n300 DP_OP_94J1_122_9915_n271 DP_OP_94J1_122_9915_n272 DP_OP_94J1_122_9915_n273 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U179 in[45] in[53] in[61] DP_OP_94J1_122_9915_n265 DP_OP_94J1_122_9915_n266 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U178 in[69] in[77] in[85] DP_OP_94J1_122_9915_n263 DP_OP_94J1_122_9915_n264 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U177 in[93] in[101] in[109] DP_OP_94J1_122_9915_n261 DP_OP_94J1_122_9915_n262 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U174 in[9] in[65] in[17] DP_OP_94J1_122_9915_n255 DP_OP_94J1_122_9915_n256 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U171 in[57] in[41] in[49] DP_OP_94J1_122_9915_n249 DP_OP_94J1_122_9915_n250 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U169 DP_OP_94J1_122_9915_n299 DP_OP_94J1_122_9915_n246 DP_OP_94J1_122_9915_n297 DP_OP_94J1_122_9915_n247 DP_OP_94J1_122_9915_n248 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U166 DP_OP_94J1_122_9915_n285 DP_OP_94J1_122_9915_n281 DP_OP_94J1_122_9915_n287 DP_OP_94J1_122_9915_n241 DP_OP_94J1_122_9915_n242 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U165 DP_OP_94J1_122_9915_n289 DP_OP_94J1_122_9915_n291 DP_OP_94J1_122_9915_n293 DP_OP_94J1_122_9915_n239 DP_OP_94J1_122_9915_n240 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U163 DP_OP_94J1_122_9915_n258 n215 DP_OP_94J1_122_9915_n256 DP_OP_94J1_122_9915_n235 DP_OP_94J1_122_9915_n236 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U162 DP_OP_94J1_122_9915_n266 DP_OP_94J1_122_9915_n254 DP_OP_94J1_122_9915_n264 DP_OP_94J1_122_9915_n233 DP_OP_94J1_122_9915_n234 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U156 DP_OP_94J1_122_9915_n234 DP_OP_94J1_122_9915_n236 n100 DP_OP_94J1_122_9915_n224 DP_OP_94J1_122_9915_n225 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U148 in[2] in[106] in[10] DP_OP_94J1_122_9915_n211 DP_OP_94J1_122_9915_n212 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U146 in[86] in[26] in[34] DP_OP_94J1_122_9915_n207 DP_OP_94J1_122_9915_n208 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U143 in[126] in[50] in[114] DP_OP_94J1_122_9915_n201 DP_OP_94J1_122_9915_n202 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U142 in[58] in[90] in[66] DP_OP_94J1_122_9915_n199 DP_OP_94J1_122_9915_n200 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U141 in[98] in[74] in[82] DP_OP_94J1_122_9915_n197 DP_OP_94J1_122_9915_n198 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U139 DP_OP_94J1_122_9915_n267 DP_OP_94J1_122_9915_n194 DP_OP_94J1_122_9915_n265 DP_OP_94J1_122_9915_n195 DP_OP_94J1_122_9915_n196 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U137 DP_OP_94J1_122_9915_n263 DP_OP_94J1_122_9915_n249 DP_OP_94J1_122_9915_n191 DP_OP_94J1_122_9915_n192 DP_OP_94J1_122_9915_n193 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U136 DP_OP_94J1_122_9915_n251 DP_OP_94J1_122_9915_n257 DP_OP_94J1_122_9915_n261 DP_OP_94J1_122_9915_n189 DP_OP_94J1_122_9915_n190 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U135 DP_OP_94J1_122_9915_n253 DP_OP_94J1_122_9915_n259 DP_OP_94J1_122_9915_n255 DP_OP_94J1_122_9915_n187 DP_OP_94J1_122_9915_n188 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U133 DP_OP_94J1_122_9915_n247 DP_OP_94J1_122_9915_n241 n168 DP_OP_94J1_122_9915_n185 DP_OP_94J1_122_9915_n186 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U131 DP_OP_94J1_122_9915_n210 DP_OP_94J1_122_9915_n202 n31 DP_OP_94J1_122_9915_n182 DP_OP_94J1_122_9915_n183 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U130 DP_OP_94J1_122_9915_n214 DP_OP_94J1_122_9915_n204 DP_OP_94J1_122_9915_n216 DP_OP_94J1_122_9915_n179 DP_OP_94J1_122_9915_n180 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U125 DP_OP_94J1_122_9915_n237 DP_OP_94J1_122_9915_n235 DP_OP_94J1_122_9915_n233 DP_OP_94J1_122_9915_n170 DP_OP_94J1_122_9915_n171 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U123 DP_OP_94J1_122_9915_n228 DP_OP_94J1_122_9915_n231 DP_OP_94J1_122_9915_n167 DP_OP_94J1_122_9915_n168 DP_OP_94J1_122_9915_n169 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U113 in[47] in[115] in[55] DP_OP_94J1_122_9915_n151 DP_OP_94J1_122_9915_n152 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U112 in[63] in[3] in[71] DP_OP_94J1_122_9915_n149 DP_OP_94J1_122_9915_n150 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U111 in[79] in[99] in[11] DP_OP_94J1_122_9915_n147 DP_OP_94J1_122_9915_n148 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U109 in[95] in[27] in[103] DP_OP_94J1_122_9915_n143 DP_OP_94J1_122_9915_n144 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U106 in[91] in[51] in[83] DP_OP_94J1_122_9915_n137 DP_OP_94J1_122_9915_n138 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U105 in[75] in[59] in[67] DP_OP_94J1_122_9915_n135 DP_OP_94J1_122_9915_n136 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U101 DP_OP_94J1_122_9915_n211 DP_OP_94J1_122_9915_n129 DP_OP_94J1_122_9915_n197 DP_OP_94J1_122_9915_n130 DP_OP_94J1_122_9915_n131 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U100 DP_OP_94J1_122_9915_n209 n48 DP_OP_94J1_122_9915_n199 DP_OP_94J1_122_9915_n127 DP_OP_94J1_122_9915_n128 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U99 DP_OP_94J1_122_9915_n207 DP_OP_94J1_122_9915_n203 DP_OP_94J1_122_9915_n201 DP_OP_94J1_122_9915_n125 DP_OP_94J1_122_9915_n126 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U93 DP_OP_94J1_122_9915_n152 DP_OP_94J1_122_9915_n154 DP_OP_94J1_122_9915_n144 DP_OP_94J1_122_9915_n115 DP_OP_94J1_122_9915_n116 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U89 n157 DP_OP_94J1_122_9915_n179 DP_OP_94J1_122_9915_n182 DP_OP_94J1_122_9915_n110 DP_OP_94J1_122_9915_n111 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U84 DP_OP_94J1_122_9915_n124 n167 DP_OP_94J1_122_9915_n170 DP_OP_94J1_122_9915_n102 DP_OP_94J1_122_9915_n103 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U82 DP_OP_94J1_122_9915_n172 DP_OP_94J1_122_9915_n114 n101 DP_OP_94J1_122_9915_n99 DP_OP_94J1_122_9915_n100 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U68 DP_OP_94J1_122_9915_n147 DP_OP_94J1_122_9915_n143 DP_OP_94J1_122_9915_n135 DP_OP_94J1_122_9915_n78 DP_OP_94J1_122_9915_n79 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U66 DP_OP_94J1_122_9915_n125 DP_OP_94J1_122_9915_n133 DP_OP_94J1_122_9915_n130 DP_OP_94J1_122_9915_n74 DP_OP_94J1_122_9915_n75 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U62 DP_OP_94J1_122_9915_n81 DP_OP_94J1_122_9915_n117 DP_OP_94J1_122_9915_n79 DP_OP_94J1_122_9915_n67 DP_OP_94J1_122_9915_n68 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U61 DP_OP_94J1_122_9915_n75 DP_OP_94J1_122_9915_n113 DP_OP_94J1_122_9915_n107 DP_OP_94J1_122_9915_n65 DP_OP_94J1_122_9915_n66 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U58 DP_OP_94J1_122_9915_n71 DP_OP_94J1_122_9915_n68 n30 DP_OP_94J1_122_9915_n61 DP_OP_94J1_122_9915_n62 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U53 DP_OP_94J1_122_9915_n76 DP_OP_94J1_122_9915_n83 DP_OP_94J1_122_9915_n80 DP_OP_94J1_122_9915_n51 DP_OP_94J1_122_9915_n52 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U50 DP_OP_94J1_122_9915_n67 DP_OP_94J1_122_9915_n52 DP_OP_94J1_122_9915_n70 DP_OP_94J1_122_9915_n46 DP_OP_94J1_122_9915_n47 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U49 DP_OP_94J1_122_9915_n50 DP_OP_94J1_122_9915_n65 DP_OP_94J1_122_9915_n63 DP_OP_94J1_122_9915_n44 DP_OP_94J1_122_9915_n45 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U44 DP_OP_94J1_122_9915_n46 DP_OP_94J1_122_9915_n49 n160 DP_OP_94J1_122_9915_n37 DP_OP_94J1_122_9915_n38 FAx1_ASAP7_75t_R
XU3 DP_OP_94J1_122_9915_n37 n96 n197 XNOR2xp5_ASAP7_75t_R
XU4 n129 n130 DP_OP_94J1_122_9915_n91 XOR2xp5_ASAP7_75t_R
XU5 n147 DP_OP_94J1_122_9915_n227 n109 XNOR2xp5_ASAP7_75t_R
XU6 n17 n153 n136 XOR2xp5_ASAP7_75t_R
XU7 DP_OP_94J1_122_9915_n103 DP_OP_94J1_122_9915_n100 n130 XNOR2xp5_ASAP7_75t_R
XU8 n174 n175 n108 XNOR2xp5_ASAP7_75t_R
XU9 n91 n131 n90 XOR2xp5_ASAP7_75t_R
XU10 n134 n65 n84 XNOR2xp5_ASAP7_75t_R
XU11 n174 n175 n104 XOR2xp5_ASAP7_75t_R
XU12 n193 n116 INVx1_ASAP7_75t_R
XU13 n45 n91 INVx2_ASAP7_75t_R
XU14 n57 n56 n44 XNOR2xp5_ASAP7_75t_R
XU15 n154 n30 INVx2_ASAP7_75t_R
XU16 DP_OP_94J1_122_9915_n123 n183 DP_OP_94J1_122_9915_n71 XOR2xp5_ASAP7_75t_R
XU17 n176 n156 DP_OP_94J1_122_9915_n176 XNOR2xp5_ASAP7_75t_R
XU18 n71 n70 DP_OP_94J1_122_9915_n227 XNOR2xp5_ASAP7_75t_R
XU19 DP_OP_94J1_122_9915_n131 n16 n64 XNOR2xp5_ASAP7_75t_R
XU20 n15 n37 n176 XNOR2xp5_ASAP7_75t_R
XU21 n141 n140 n101 XNOR2xp5_ASAP7_75t_R
XU22 in[7] in[15] DP_OP_94J1_122_9915_n129 XNOR2xp5_ASAP7_75t_R
XU23 in[81] n88 n87 XNOR2xp5_ASAP7_75t_R
XU24 in[117] in[1] n88 XOR2xp5_ASAP7_75t_R
XU25 in[123] in[43] n139 XOR2xp5_ASAP7_75t_R
XU26 DP_OP_94J1_122_9915_n198 n168 INVx1_ASAP7_75t_R
XU27 n5 TIEHIx1_ASAP7_75t_R
XU28 n5 out[9] INVx1_ASAP7_75t_R
XU29 n5 out[10] INVx1_ASAP7_75t_R
XU30 n5 out[11] INVx1_ASAP7_75t_R
XU31 n5 out[12] INVx1_ASAP7_75t_R
XU32 DP_OP_94J1_122_9915_n195 n6 DP_OP_94J1_122_9915_n124 XOR2xp5_ASAP7_75t_R
XU33 n103 DP_OP_94J1_122_9915_n189 n6 XNOR2xp5_ASAP7_75t_R
XU34 n63 n197 n32 n127 NAND3xp33_ASAP7_75t_R
XU35 n51 n136 DP_OP_94J1_122_9915_n40 XNOR2xp5_ASAP7_75t_R
XU36 DP_OP_94J1_122_9915_n102 n154 BUFx2_ASAP7_75t_R
XU37 DP_OP_94J1_122_9915_n195 n103 DP_OP_94J1_122_9915_n189 n7 MAJIxp5_ASAP7_75t_R
XU38 DP_OP_94J1_122_9915_n195 n103 DP_OP_94J1_122_9915_n189 DP_OP_94J1_122_9915_n123 MAJx2_ASAP7_75t_R
XU39 n8 DP_OP_94J1_122_9915_n248 n100 XOR2x2_ASAP7_75t_R
XU40 DP_OP_94J1_122_9915_n279 n47 n8 XOR2xp5_ASAP7_75t_R
XU41 n55 n54 n32 AND2x2_ASAP7_75t_R
XU42 in[14] in[6] DP_OP_94J1_122_9915_n132 NAND2xp5_ASAP7_75t_R
XU43 n46 n123 n122 NAND2xp5_ASAP7_75t_R
XU44 DP_OP_94J1_122_9915_n207 DP_OP_94J1_122_9915_n203 DP_OP_94J1_122_9915_n201 n9 MAJIxp5_ASAP7_75t_R
XU45 n13 n29 n66 n10 MAJIxp5_ASAP7_75t_R
XU46 n13 n29 n66 n11 MAJIxp5_ASAP7_75t_R
XU47 DP_OP_94J1_122_9915_n200 DP_OP_94J1_122_9915_n206 DP_OP_94J1_122_9915_n212 n12 MAJIxp5_ASAP7_75t_R
XU48 n129 n130 n13 XNOR2xp5_ASAP7_75t_R
XU49 DP_OP_94J1_122_9915_n37 n96 n14 XOR2xp5_ASAP7_75t_R
XU50 n34 DP_OP_94J1_122_9915_n283 DP_OP_94J1_122_9915_n295 n15 MAJIxp5_ASAP7_75t_R
XU51 n34 DP_OP_94J1_122_9915_n283 DP_OP_94J1_122_9915_n295 DP_OP_94J1_122_9915_n244 MAJx2_ASAP7_75t_R
XU52 DP_OP_94J1_122_9915_n200 DP_OP_94J1_122_9915_n206 DP_OP_94J1_122_9915_n212 n16 MAJx2_ASAP7_75t_R
XU53 DP_OP_94J1_122_9915_n47 DP_OP_94J1_122_9915_n61 n17 XNOR2xp5_ASAP7_75t_R
XU54 in[4] in[28] in[36] n18 MAJIxp5_ASAP7_75t_R
XU55 n196 n98 n19 XOR2xp5_ASAP7_75t_R
XU56 n196 n98 n59 XOR2xp5_ASAP7_75t_R
XU57 DP_OP_94J1_122_9915_n226 DP_OP_94J1_122_9915_n176 n131 XOR2x2_ASAP7_75t_R
XU58 n84 n193 n196 XNOR2x2_ASAP7_75t_R
XU59 DP_OP_94J1_122_9915_n99 n118 BUFx4_ASAP7_75t_R
XU60 DP_OP_94J1_122_9915_n168 n111 BUFx4_ASAP7_75t_R
XU61 DP_OP_94J1_122_9915_n240 n25 BUFx4_ASAP7_75t_R
XU62 in[30] in[38] in[22] n20 MAJIxp5_ASAP7_75t_R
XU63 in[13] in[5] n21 XOR2xp5_ASAP7_75t_R
XU64 n57 n56 n22 XOR2xp5_ASAP7_75t_R
XU65 n60 n19 n23 XOR2xp5_ASAP7_75t_R
XU66 DP_OP_94J1_122_9915_n245 n172 n24 XOR2xp5_ASAP7_75t_R
XU67 in[81] n88 n26 XOR2xp5_ASAP7_75t_R
XU68 n131 n45 n27 XNOR2xp5_ASAP7_75t_R
XU69 n71 n70 n28 XOR2xp5_ASAP7_75t_R
XU70 DP_OP_94J1_122_9915_n239 n159 BUFx4_ASAP7_75t_R
XU71 n39 n73 INVx3_ASAP7_75t_R
XU72 n78 DP_OP_94J1_122_9915_n161 n206 n29 MAJx2_ASAP7_75t_R
XU73 n159 n31 INVx3_ASAP7_75t_R
XU74 DP_OP_94J1_122_9915_n171 n45 BUFx4_ASAP7_75t_R
XU75 in[13] in[5] n34 XNOR2xp5_ASAP7_75t_R
XU76 n45 n131 n35 XOR2x2_ASAP7_75t_R
XU77 DP_OP_94J1_122_9915_n183 n36 HB1xp67_ASAP7_75t_R
XU78 n43 n170 HB1xp67_ASAP7_75t_R
XU79 n170 n37 INVx1_ASAP7_75t_R
XU80 n50 n163 n38 OR2x2_ASAP7_75t_R
XU81 n37 n15 n102 NOR2xp33_ASAP7_75t_R
XU82 n75 n39 BUFx6f_ASAP7_75t_R
XU83 DP_OP_94J1_122_9915_n110 n76 n75 XNOR2x2_ASAP7_75t_R
XU84 n78 n206 DP_OP_94J1_122_9915_n161 n40 MAJIxp5_ASAP7_75t_R
XU85 DP_OP_94J1_122_9915_n245 n172 n41 XNOR2xp5_ASAP7_75t_R
XU86 n60 n59 n42 XNOR2xp5_ASAP7_75t_R
XU87 in[86] in[26] in[34] n43 FAx1_ASAP7_75t_R
XU88 n171 DP_OP_94J1_122_9915_n57 n42 n46 MAJIxp5_ASAP7_75t_R
XU89 n121 n123 n63 NAND2xp33_ASAP7_75t_R
XU90 DP_OP_94J1_122_9915_n244 DP_OP_94J1_122_9915_n208 n72 NOR2xp33_ASAP7_75t_R
XU91 DP_OP_94J1_122_9915_n276 DP_OP_94J1_122_9915_n274 n69 NAND2xp33_ASAP7_75t_R
XU92 in[13] in[5] DP_OP_94J1_122_9915_n194 NAND2xp5_ASAP7_75t_R
XU93 n69 n71 n68 NAND2xp33_ASAP7_75t_R
XU94 in[7] in[15] n213 NAND2xp33_ASAP7_75t_R
XU95 DP_OP_94J1_122_9915_n77 DP_OP_94J1_122_9915_n120 n183 XNOR2xp5_ASAP7_75t_R
XU96 in[21] n62 n47 XOR2xp5_ASAP7_75t_R
XU97 in[122] in[102] in[94] n48 MAJIxp5_ASAP7_75t_R
XU98 DP_OP_94J1_122_9915_n276 DP_OP_94J1_122_9915_n274 n49 OR2x2_ASAP7_75t_R
XU99 DP_OP_94J1_122_9915_n56 DP_OP_94J1_122_9915_n45 n136 n50 MAJIxp5_ASAP7_75t_R
XU100 in[127] n139 n103 XOR2xp5_ASAP7_75t_R
XU101 n14 n38 n126 AND2x2_ASAP7_75t_R
XU102 n111 n155 INVx2_ASAP7_75t_R
XU103 n118 n134 INVx2_ASAP7_75t_R
XU104 n162 n161 INVx2_ASAP7_75t_R
XU105 n117 n65 INVxp67_ASAP7_75t_R
XU106 n102 n135 n57 NOR2xp67_ASAP7_75t_R
XU107 n72 n115 n135 NOR2xp33_ASAP7_75t_R
XU108 DP_OP_94J1_122_9915_n196 n156 INVxp67_ASAP7_75t_R
XU109 n25 n173 INVx2_ASAP7_75t_R
XU110 DP_OP_94J1_122_9915_n200 n177 DP_OP_94J1_122_9915_n178 XOR2xp5_ASAP7_75t_R
XU111 in[38] in[30] n133 XOR2xp5_ASAP7_75t_R
XU112 n210 DP_OP_94J1_122_9915_n40 n123 OR2x2_ASAP7_75t_R
XU113 n116 DP_OP_94J1_122_9915_n66 n118 n153 MAJx2_ASAP7_75t_R
XU114 DP_OP_94J1_122_9915_n56 n52 n51 XNOR2xp5_ASAP7_75t_R
XU115 n114 n52 INVxp67_ASAP7_75t_R
XU116 DP_OP_94J1_122_9915_n62 n53 n73 DP_OP_94J1_122_9915_n56 MAJIxp5_ASAP7_75t_R
XU117 n125 n127 n158 out[7] NAND3xp33_ASAP7_75t_R
XU118 n53 n39 n74 XNOR2xp5_ASAP7_75t_R
XU119 DP_OP_94J1_122_9915_n162 n44 n216 n53 MAJIxp5_ASAP7_75t_R
XU120 n163 n50 n54 NAND2xp5_ASAP7_75t_R
XU121 n210 DP_OP_94J1_122_9915_n40 n55 NAND2xp5_ASAP7_75t_R
XU122 DP_OP_94J1_122_9915_n116 DP_OP_94J1_122_9915_n126 n57 DP_OP_94J1_122_9915_n105 MAJIxp5_ASAP7_75t_R
XU123 DP_OP_94J1_122_9915_n126 DP_OP_94J1_122_9915_n116 n56 XOR2xp5_ASAP7_75t_R
XU124 DP_OP_94J1_122_9915_n193 DP_OP_94J1_122_9915_n188 DP_OP_94J1_122_9915_n190 DP_OP_94J1_122_9915_n172 MAJIxp5_ASAP7_75t_R
XU125 DP_OP_94J1_122_9915_n193 n58 DP_OP_94J1_122_9915_n173 XOR2xp5_ASAP7_75t_R
XU126 DP_OP_94J1_122_9915_n188 DP_OP_94J1_122_9915_n190 n58 XNOR2xp5_ASAP7_75t_R
XU127 n13 n29 n66 n171 MAJIxp5_ASAP7_75t_R
XU128 n195 n61 n66 XNOR2xp5_ASAP7_75t_R
XU129 n10 DP_OP_94J1_122_9915_n57 n42 n121 MAJIxp5_ASAP7_75t_R
XU130 n194 n195 n108 n60 MAJIxp5_ASAP7_75t_R
XU131 n104 n194 n61 XOR2xp5_ASAP7_75t_R
XU132 in[21] in[37] in[29] DP_OP_94J1_122_9915_n267 MAJIxp5_ASAP7_75t_R
XU133 in[37] in[29] n62 XOR2xp5_ASAP7_75t_R
XU134 DP_OP_94J1_122_9915_n128 DP_OP_94J1_122_9915_n131 n12 DP_OP_94J1_122_9915_n107 MAJIxp5_ASAP7_75t_R
XU135 DP_OP_94J1_122_9915_n128 n64 DP_OP_94J1_122_9915_n108 XNOR2xp5_ASAP7_75t_R
XU136 n66 DP_OP_94J1_122_9915_n91 n208 XNOR2xp5_ASAP7_75t_R
XU137 n67 n27 n78 XNOR2xp5_ASAP7_75t_R
XU138 n35 n67 n205 XNOR2xp5_ASAP7_75t_R
XU139 DP_OP_94J1_122_9915_n169 DP_OP_94J1_122_9915_n221 n67 XNOR2xp5_ASAP7_75t_R
XU140 n49 n68 DP_OP_94J1_122_9915_n226 NAND2xp5_ASAP7_75t_R
XU141 DP_OP_94J1_122_9915_n274 DP_OP_94J1_122_9915_n276 n70 XNOR2xp5_ASAP7_75t_R
XU142 n81 n26 n71 XOR2xp5_ASAP7_75t_R
XU143 n74 DP_OP_94J1_122_9915_n62 DP_OP_94J1_122_9915_n57 XNOR2xp5_ASAP7_75t_R
XU144 DP_OP_94J1_122_9915_n73 DP_OP_94J1_122_9915_n105 n76 XNOR2xp5_ASAP7_75t_R
XU145 n45 DP_OP_94J1_122_9915_n226 DP_OP_94J1_122_9915_n176 DP_OP_94J1_122_9915_n162 MAJx2_ASAP7_75t_R
XU146 n77 DP_OP_94J1_122_9915_n225 n204 n206 MAJIxp5_ASAP7_75t_R
XU147 n147 n28 n77 XNOR2xp5_ASAP7_75t_R
XU148 n24 n107 n147 XNOR2xp5_ASAP7_75t_R
XU149 n107 n41 DP_OP_94J1_122_9915_n227 DP_OP_94J1_122_9915_n221 MAJIxp5_ASAP7_75t_R
XU150 n80 n79 DP_OP_94J1_122_9915_n50 XNOR2xp5_ASAP7_75t_R
XU151 n166 DP_OP_94J1_122_9915_n74 n79 XOR2xp5_ASAP7_75t_R
XU152 n166 n80 DP_OP_94J1_122_9915_n74 DP_OP_94J1_122_9915_n49 MAJIxp5_ASAP7_75t_R
XU153 DP_OP_94J1_122_9915_n115 DP_OP_94J1_122_9915_n84 DP_OP_94J1_122_9915_n127 n80 MAJIxp5_ASAP7_75t_R
XU154 DP_OP_94J1_122_9915_n250 DP_OP_94J1_122_9915_n262 n81 XNOR2xp5_ASAP7_75t_R
XU155 n20 DP_OP_94J1_122_9915_n213 DP_OP_94J1_122_9915_n132 DP_OP_94J1_122_9915_n133 MAJIxp5_ASAP7_75t_R
XU156 n83 n82 DP_OP_94J1_122_9915_n134 XNOR2xp5_ASAP7_75t_R
XU157 DP_OP_94J1_122_9915_n132 DP_OP_94J1_122_9915_n213 n82 XNOR2xp5_ASAP7_75t_R
XU158 in[30] in[38] in[22] n83 MAJx2_ASAP7_75t_R
XU159 n120 n119 n163 XNOR2xp5_ASAP7_75t_R
XU160 n179 n85 n178 NAND2xp33_ASAP7_75t_R
XU161 n126 n85 n125 NAND2xp5_ASAP7_75t_R
XU162 n122 n32 n85 NAND2xp5_ASAP7_75t_R
XU163 n86 n21 DP_OP_94J1_122_9915_n245 XNOR2xp5_ASAP7_75t_R
XU164 DP_OP_94J1_122_9915_n283 DP_OP_94J1_122_9915_n295 n86 XNOR2xp5_ASAP7_75t_R
XU165 DP_OP_94J1_122_9915_n262 n87 DP_OP_94J1_122_9915_n250 DP_OP_94J1_122_9915_n237 MAJIxp5_ASAP7_75t_R
XU166 DP_OP_94J1_122_9915_n162 n89 n194 XNOR2xp5_ASAP7_75t_R
XU167 n216 n22 n89 XNOR2xp5_ASAP7_75t_R
XU168 DP_OP_94J1_122_9915_n169 n90 DP_OP_94J1_122_9915_n221 n195 MAJx2_ASAP7_75t_R
XU169 n212 n92 out[6] XOR2xp5_ASAP7_75t_R
XU170 DP_OP_94J1_122_9915_n40 n210 n121 n92 MAJIxp5_ASAP7_75t_R
XU171 n9 DP_OP_94J1_122_9915_n133 DP_OP_94J1_122_9915_n130 n93 FAx1_ASAP7_75t_R
XU172 in[45] in[53] in[61] n94 MAJIxp5_ASAP7_75t_R
XU173 n97 DP_OP_94J1_122_9915_n37 n180 NAND2xp33_ASAP7_75t_R
XU174 in[78] in[18] n192 XOR2xp5_ASAP7_75t_R
XU175 in[102] in[122] n201 XOR2xp5_ASAP7_75t_R
XU176 in[16] in[8] n198 XOR2xp5_ASAP7_75t_R
XU177 DP_OP_94J1_122_9915_n37 n97 n164 OR2x2_ASAP7_75t_R
XU178 n129 DP_OP_94J1_122_9915_n103 DP_OP_94J1_122_9915_n100 n95 MAJIxp5_ASAP7_75t_R
XU179 n120 DP_OP_94J1_122_9915_n44 DP_OP_94J1_122_9915_n38 n96 MAJIxp5_ASAP7_75t_R
XU180 n111 DP_OP_94J1_122_9915_n108 n174 XOR2x2_ASAP7_75t_R
XU181 n155 DP_OP_94J1_122_9915_n108 n151 n193 MAJx3_ASAP7_75t_R
XU182 n120 DP_OP_94J1_122_9915_n44 DP_OP_94J1_122_9915_n38 n97 MAJx2_ASAP7_75t_R
XU183 n129 DP_OP_94J1_122_9915_n103 DP_OP_94J1_122_9915_n100 n98 MAJx2_ASAP7_75t_R
XU184 DP_OP_94J1_122_9915_n187 n105 BUFx4_ASAP7_75t_R
XU185 DP_OP_94J1_122_9915_n272 n148 BUFx4_ASAP7_75t_R
XU186 in[35] in[119] in[111] n99 MAJIxp5_ASAP7_75t_R
XU187 DP_OP_94J1_122_9915_n136 DP_OP_94J1_122_9915_n150 n140 XNOR2x2_ASAP7_75t_R
XU188 in[63] in[3] in[71] n110 MAJx2_ASAP7_75t_R
XU189 DP_OP_94J1_122_9915_n209 n48 DP_OP_94J1_122_9915_n199 n113 MAJx2_ASAP7_75t_R
XU190 n105 n141 INVx3_ASAP7_75t_R
XU191 DP_OP_94J1_122_9915_n280 n106 HB1xp67_ASAP7_75t_R
XU192 n148 n107 INVx3_ASAP7_75t_R
XU193 n18 DP_OP_94J1_122_9915_n246 DP_OP_94J1_122_9915_n297 n112 FAx1_ASAP7_75t_R
XU194 DP_OP_94J1_122_9915_n50 DP_OP_94J1_122_9915_n65 DP_OP_94J1_122_9915_n63 n114 FAx1_ASAP7_75t_R
XU195 DP_OP_94J1_122_9915_n267 DP_OP_94J1_122_9915_n194 n94 n115 FAx1_ASAP7_75t_R
XU196 n93 DP_OP_94J1_122_9915_n113 DP_OP_94J1_122_9915_n107 n117 FAx1_ASAP7_75t_R
XU197 n112 n47 DP_OP_94J1_122_9915_n279 DP_OP_94J1_122_9915_n231 MAJIxp5_ASAP7_75t_R
XU198 DP_OP_94J1_122_9915_n44 DP_OP_94J1_122_9915_n38 n119 XOR2xp5_ASAP7_75t_R
XU199 n153 DP_OP_94J1_122_9915_n47 DP_OP_94J1_122_9915_n61 n120 MAJIxp5_ASAP7_75t_R
XU200 in[64] in[48] in[56] DP_OP_94J1_122_9915_n285 MAJIxp5_ASAP7_75t_R
XU201 in[64] n124 DP_OP_94J1_122_9915_n286 XNOR2xp5_ASAP7_75t_R
XU202 in[48] in[56] n124 XOR2xp5_ASAP7_75t_R
XU203 in[46] in[62] in[54] DP_OP_94J1_122_9915_n213 MAJIxp5_ASAP7_75t_R
XU204 in[46] n128 DP_OP_94J1_122_9915_n214 XNOR2xp5_ASAP7_75t_R
XU205 in[62] in[54] n128 XOR2xp5_ASAP7_75t_R
XU206 DP_OP_94J1_122_9915_n224 DP_OP_94J1_122_9915_n173 n186 n129 MAJIxp5_ASAP7_75t_R
XU207 DP_OP_94J1_122_9915_n273 DP_OP_94J1_122_9915_n275 DP_OP_94J1_122_9915_n277 n204 MAJIxp5_ASAP7_75t_R
XU208 in[113] in[25] in[97] DP_OP_94J1_122_9915_n253 MAJIxp5_ASAP7_75t_R
XU209 in[113] n132 DP_OP_94J1_122_9915_n254 XNOR2xp5_ASAP7_75t_R
XU210 in[25] in[97] n132 XOR2xp5_ASAP7_75t_R
XU211 in[22] n133 DP_OP_94J1_122_9915_n216 XNOR2xp5_ASAP7_75t_R
XU212 n99 DP_OP_94J1_122_9915_n139 DP_OP_94J1_122_9915_n145 DP_OP_94J1_122_9915_n76 MAJIxp5_ASAP7_75t_R
XU213 n138 n137 DP_OP_94J1_122_9915_n77 XNOR2xp5_ASAP7_75t_R
XU214 DP_OP_94J1_122_9915_n139 DP_OP_94J1_122_9915_n145 n137 XNOR2xp5_ASAP7_75t_R
XU215 in[35] in[119] in[111] n138 MAJx2_ASAP7_75t_R
XU216 in[127] in[123] in[43] DP_OP_94J1_122_9915_n139 MAJIxp5_ASAP7_75t_R
XU217 n141 DP_OP_94J1_122_9915_n136 DP_OP_94J1_122_9915_n150 DP_OP_94J1_122_9915_n120 MAJIxp5_ASAP7_75t_R
XU218 DP_OP_94J1_122_9915_n149 DP_OP_94J1_122_9915_n137 DP_OP_94J1_122_9915_n151 DP_OP_94J1_122_9915_n80 MAJIxp5_ASAP7_75t_R
XU219 n110 n142 DP_OP_94J1_122_9915_n81 XNOR2xp5_ASAP7_75t_R
XU220 DP_OP_94J1_122_9915_n137 DP_OP_94J1_122_9915_n151 n142 XNOR2xp5_ASAP7_75t_R
XU221 in[23] in[39] in[31] DP_OP_94J1_122_9915_n153 MAJIxp5_ASAP7_75t_R
XU222 in[23] n143 DP_OP_94J1_122_9915_n154 XNOR2xp5_ASAP7_75t_R
XU223 in[39] in[31] n143 XOR2xp5_ASAP7_75t_R
XU224 n144 DP_OP_94J1_122_9915_n115 DP_OP_94J1_122_9915_n73 XNOR2xp5_ASAP7_75t_R
XU225 n113 DP_OP_94J1_122_9915_n84 n144 XNOR2xp5_ASAP7_75t_R
XU226 in[19] in[87] in[107] DP_OP_94J1_122_9915_n145 MAJIxp5_ASAP7_75t_R
XU227 in[19] n145 DP_OP_94J1_122_9915_n146 XNOR2xp5_ASAP7_75t_R
XU228 in[87] in[107] n145 XOR2xp5_ASAP7_75t_R
XU229 in[125] in[121] in[89] DP_OP_94J1_122_9915_n257 MAJIxp5_ASAP7_75t_R
XU230 in[125] n146 DP_OP_94J1_122_9915_n258 XNOR2xp5_ASAP7_75t_R
XU231 in[121] in[89] n146 XOR2xp5_ASAP7_75t_R
XU232 n164 n178 out[8] NAND2xp33_ASAP7_75t_R
XU233 n194 n108 n195 n149 MAJIxp5_ASAP7_75t_R
XU234 in[58] in[90] in[66] n150 FAx1_ASAP7_75t_R
XU235 DP_OP_94J1_122_9915_n111 n151 BUFx4_ASAP7_75t_R
XU236 n150 n177 n152 XNOR2xp5_ASAP7_75t_R
XU237 n163 n50 n212 XNOR2xp5_ASAP7_75t_R
XU238 DP_OP_94J1_122_9915_n185 DP_OP_94J1_122_9915_n109 BUFx4_ASAP7_75t_R
XU239 n151 n175 INVx3_ASAP7_75t_R
XU240 DP_OP_94J1_122_9915_n109 n157 INVx3_ASAP7_75t_R
XU241 DP_OP_94J1_122_9915_n186 n162 BUFx4_ASAP7_75t_R
XU242 n106 DP_OP_94J1_122_9915_n271 INVx1_ASAP7_75t_R
XU243 n38 n180 n179 AND2x2_ASAP7_75t_R
XU244 n14 n38 n158 OR2x2_ASAP7_75t_R
XU245 DP_OP_94J1_122_9915_n51 DP_OP_94J1_122_9915_n36 BUFx4_ASAP7_75t_R
XU246 DP_OP_94J1_122_9915_n36 n160 INVx3_ASAP7_75t_R
XU247 DP_OP_94J1_122_9915_n138 n199 BUFx4_ASAP7_75t_R
XU248 n36 DP_OP_94J1_122_9915_n167 INVx1_ASAP7_75t_R
XU249 DP_OP_94J1_122_9915_n78 DP_OP_94J1_122_9915_n48 BUFx4_ASAP7_75t_R
XU250 DP_OP_94J1_122_9915_n153 n213 DP_OP_94J1_122_9915_n83 NOR2x1_ASAP7_75t_R
XU251 DP_OP_94J1_122_9915_n120 DP_OP_94J1_122_9915_n77 n165 OR2x2_ASAP7_75t_R
XU252 DP_OP_94J1_122_9915_n48 n166 INVx3_ASAP7_75t_R
XU253 DP_OP_94J1_122_9915_n146 n191 n167 XNOR2xp5_ASAP7_75t_R
XU254 n199 n169 INVx3_ASAP7_75t_R
XU255 n25 DP_OP_94J1_122_9915_n242 DP_OP_94J1_122_9915_n245 DP_OP_94J1_122_9915_n228 MAJIxp5_ASAP7_75t_R
XU256 DP_OP_94J1_122_9915_n242 n173 n172 XNOR2xp5_ASAP7_75t_R
XU257 n210 DP_OP_94J1_122_9915_n40 n211 XNOR2xp5_ASAP7_75t_R
XU258 DP_OP_94J1_122_9915_n206 DP_OP_94J1_122_9915_n212 n177 XNOR2xp5_ASAP7_75t_R
XU259 n181 n165 DP_OP_94J1_122_9915_n70 NAND2xp5_ASAP7_75t_R
XU260 n7 n182 n181 NAND2xp33_ASAP7_75t_R
XU261 DP_OP_94J1_122_9915_n77 DP_OP_94J1_122_9915_n120 n182 NAND2xp5_ASAP7_75t_R
XU262 in[111] n184 DP_OP_94J1_122_9915_n142 XNOR2xp5_ASAP7_75t_R
XU263 in[119] in[35] n184 XOR2xp5_ASAP7_75t_R
XU264 DP_OP_94J1_122_9915_n224 n185 DP_OP_94J1_122_9915_n161 XNOR2xp5_ASAP7_75t_R
XU265 n186 DP_OP_94J1_122_9915_n173 n185 XOR2xp5_ASAP7_75t_R
XU266 n187 n162 n186 XNOR2xp5_ASAP7_75t_R
XU267 DP_OP_94J1_122_9915_n180 n152 n187 XOR2xp5_ASAP7_75t_R
XU268 in[112] in[96] in[104] DP_OP_94J1_122_9915_n289 MAJIxp5_ASAP7_75t_R
XU269 in[112] n188 DP_OP_94J1_122_9915_n290 XNOR2xp5_ASAP7_75t_R
XU270 in[96] in[104] n188 XOR2xp5_ASAP7_75t_R
XU271 DP_OP_94J1_122_9915_n110 DP_OP_94J1_122_9915_n73 DP_OP_94J1_122_9915_n105 DP_OP_94J1_122_9915_n63 MAJIxp5_ASAP7_75t_R
XU272 in[110] in[118] in[42] DP_OP_94J1_122_9915_n203 MAJIxp5_ASAP7_75t_R
XU273 in[110] n189 DP_OP_94J1_122_9915_n204 XNOR2xp5_ASAP7_75t_R
XU274 in[118] in[42] n189 XOR2xp5_ASAP7_75t_R
XU275 in[116] in[120] in[124] DP_OP_94J1_122_9915_n291 MAJIxp5_ASAP7_75t_R
XU276 in[116] n190 DP_OP_94J1_122_9915_n292 XNOR2xp5_ASAP7_75t_R
XU277 in[120] in[124] n190 XOR2xp5_ASAP7_75t_R
XU278 DP_OP_94J1_122_9915_n146 DP_OP_94J1_122_9915_n142 DP_OP_94J1_122_9915_n148 DP_OP_94J1_122_9915_n117 MAJIxp5_ASAP7_75t_R
XU279 DP_OP_94J1_122_9915_n142 DP_OP_94J1_122_9915_n148 n191 XNOR2xp5_ASAP7_75t_R
XU280 in[70] in[78] in[18] DP_OP_94J1_122_9915_n209 MAJIxp5_ASAP7_75t_R
XU281 in[70] n192 DP_OP_94J1_122_9915_n210 XNOR2xp5_ASAP7_75t_R
XU282 in[20] in[12] DP_OP_94J1_122_9915_n246 NAND2xp5_ASAP7_75t_R
XU283 n161 DP_OP_94J1_122_9915_n178 DP_OP_94J1_122_9915_n180 n216 MAJIxp5_ASAP7_75t_R
XU284 n196 n95 n149 n210 MAJIxp5_ASAP7_75t_R
XU285 in[105] in[73] in[33] DP_OP_94J1_122_9915_n251 MAJIxp5_ASAP7_75t_R
XU286 in[24] in[16] in[8] DP_OP_94J1_122_9915_n281 MAJIxp5_ASAP7_75t_R
XU287 in[24] n198 DP_OP_94J1_122_9915_n282 XNOR2xp5_ASAP7_75t_R
XU288 n169 DP_OP_94J1_122_9915_n192 DP_OP_94J1_122_9915_n134 DP_OP_94J1_122_9915_n113 MAJIxp5_ASAP7_75t_R
XU289 DP_OP_94J1_122_9915_n192 n169 n200 XNOR2xp5_ASAP7_75t_R
XU290 DP_OP_94J1_122_9915_n134 n200 DP_OP_94J1_122_9915_n114 XOR2xp5_ASAP7_75t_R
XU291 in[94] n201 DP_OP_94J1_122_9915_n206 XNOR2xp5_ASAP7_75t_R
XU292 in[117] in[1] in[81] DP_OP_94J1_122_9915_n259 MAJIxp5_ASAP7_75t_R
XU293 in[14] in[6] DP_OP_94J1_122_9915_n191 HAxp5_ASAP7_75t_R
XU294 in[20] in[12] DP_OP_94J1_122_9915_n278 HAxp5_ASAP7_75t_R
XU295 DP_OP_94J1_122_9915_n277 DP_OP_94J1_122_9915_n275 n202 HAxp5_ASAP7_75t_R
XU296 DP_OP_94J1_122_9915_n273 n202 out[0] HAxp5_ASAP7_75t_R
XU297 DP_OP_94J1_122_9915_n225 n109 n203 HAxp5_ASAP7_75t_R
XU298 n204 n203 out[1] HAxp5_ASAP7_75t_R
XU299 DP_OP_94J1_122_9915_n161 n205 n207 XOR2xp5_ASAP7_75t_R
XU300 n207 n206 out[2] HAxp5_ASAP7_75t_R
XU301 n208 n40 out[3] HAxp5_ASAP7_75t_R
XU302 DP_OP_94J1_122_9915_n57 n23 n209 HAxp5_ASAP7_75t_R
XU303 n209 n11 out[4] HAxp5_ASAP7_75t_R
XU304 n211 n46 out[5] HAxp5_ASAP7_75t_R
XU305 DP_OP_94J1_122_9915_n153 n213 DP_OP_94J1_122_9915_n84 XOR2xp5_ASAP7_75t_R
XU306 in[73] in[33] n214 XOR2xp5_ASAP7_75t_R
XU307 in[105] n214 n215 XNOR2xp5_ASAP7_75t_R
.ENDS


