.SUBCKT Accumulator VSS VDD  clk rst_n in_valid partial_sum[12] partial_sum[11] partial_sum[10] partial_sum[9] partial_sum[8] partial_sum[7] partial_sum[6] partial_sum[5] partial_sum[4] partial_sum[3] partial_sum[2] partial_sum[1] partial_sum[0] result[12] result[11] result[10] result[9] result[8] result[7] result[6] result[5] result[4] result[3] result[2] result[1] result[0]
Xresult_reg_12_ VSS VDD  clk N_30 n2 n28 n14 ASYNC_DFFHx1_ASAP7_75t_L
Xresult_reg_11_ VSS VDD  clk N_29 n2 n54 n13 ASYNC_DFFHx1_ASAP7_75t_L
Xresult_reg_10_ VSS VDD  clk N_28 n2 n26 n12 ASYNC_DFFHx1_ASAP7_75t_L
Xresult_reg_9_ VSS VDD   clk N_27 n2 n29 n11 ASYNC_DFFHx1_ASAP7_75t_L
Xresult_reg_8_ VSS VDD   clk N_26 n2 n53 n10 ASYNC_DFFHx1_ASAP7_75t_L
Xresult_reg_7_ VSS VDD   clk N_25 n2 n55 n9 ASYNC_DFFHx1_ASAP7_75t_L
Xresult_reg_6_ VSS VDD   clk N_24 n2 n24 n8 ASYNC_DFFHx1_ASAP7_75t_L
Xresult_reg_5_ VSS VDD   clk N_23 n2 n30 n7 ASYNC_DFFHx1_ASAP7_75t_L
Xresult_reg_4_ VSS VDD   clk N_22 n2 n15 n6 ASYNC_DFFHx1_ASAP7_75t_L
Xresult_reg_3_ VSS VDD   clk N_21 n2 n25 n5 ASYNC_DFFHx1_ASAP7_75t_L
Xresult_reg_2_ VSS VDD   clk N_20 n2 n27 n4 ASYNC_DFFHx1_ASAP7_75t_L
Xresult_reg_1_ VSS VDD   clk N_19 n2 n23 n3 ASYNC_DFFHx1_ASAP7_75t_L
Xresult_reg_0_ VSS VDD   clk N_18 n2 n56 n1 ASYNC_DFFHx1_ASAP7_75t_L
XU31 VSS VDD  n38 result[3] INVx1_ASAP7_75t_L
XU32 VSS VDD  n39 result[5] INVx1_ASAP7_75t_L
XU33 VSS VDD  n32 result[7] INVx1_ASAP7_75t_L
XU34 VSS VDD  n33 result[9] INVx1_ASAP7_75t_L
XU35 VSS VDD  n37 result[1] INVx1_ASAP7_75t_L
XU36 VSS VDD  n121 result[0] INVx2_ASAP7_75t_L
XU37 VSS VDD  partial_sum[2] n34 INVx4_ASAP7_75t_L
XU38 VSS VDD  partial_sum[4] n47 INVx4_ASAP7_75t_L
XU39 VSS VDD  partial_sum[6] n46 INVx4_ASAP7_75t_L
XU40 VSS VDD  partial_sum[8] n45 INVx4_ASAP7_75t_L
XU41 VSS VDD  partial_sum[10] n44 INVx4_ASAP7_75t_L
XU42 VSS VDD  n4 n120 BUFx3_ASAP7_75t_L
XU43 VSS VDD  n6 n119 BUFx3_ASAP7_75t_L
XU44 VSS VDD  result[0] partial_sum[1] n48 AND2x2_ASAP7_75t_L
XU45 VSS VDD  n1 n121 BUFx3_ASAP7_75t_L
XU46 VSS VDD  n11 n33 BUFx5_ASAP7_75t_L
XU47 VSS VDD  n3 n37 BUFx5_ASAP7_75t_L
XU48 VSS VDD  n5 n38 BUFx5_ASAP7_75t_L
XU49 VSS VDD  n7 n39 BUFx5_ASAP7_75t_L
XU50 VSS VDD  n9 n32 BUFx5_ASAP7_75t_L
XU51 VSS VDD  in_valid n16 INVx4_ASAP7_75t_L
XU52 VSS VDD  in_valid n17 INVx4_ASAP7_75t_L
XU53 VSS VDD  in_valid n18 INVx4_ASAP7_75t_L
XU54 VSS VDD  in_valid n19 INVx8_ASAP7_75t_L
XU55 VSS VDD  in_valid n20 INVx4_ASAP7_75t_L
XU56 VSS VDD  in_valid n21 INVx4_ASAP7_75t_L
XU57 VSS VDD  in_valid n22 INVx4_ASAP7_75t_L
XU58 VSS VDD  in_valid n49 INVx4_ASAP7_75t_L
XU59 VSS VDD  in_valid n50 INVx4_ASAP7_75t_L
XU60 VSS VDD  rst_n n23 INVx6_ASAP7_75t_L
XU61 VSS VDD  rst_n n24 INVx6_ASAP7_75t_L
XU62 VSS VDD  rst_n n25 INVx6_ASAP7_75t_L
XU63 VSS VDD  rst_n n26 INVx6_ASAP7_75t_L
XU64 VSS VDD  rst_n n27 INVx6_ASAP7_75t_L
XU65 VSS VDD  rst_n n28 INVx6_ASAP7_75t_L
XU66 VSS VDD  rst_n n29 INVx6_ASAP7_75t_L
XU67 VSS VDD  rst_n n30 INVx6_ASAP7_75t_L
XU68 VSS VDD  result[0] partial_sum[1] n62 NAND2xp33_ASAP7_75t_L
XU69 VSS VDD  n13 n31 BUFx3_ASAP7_75t_L
XU70 VSS VDD  partial_sum[2] n63 INVx6_ASAP7_75t_L
XU71 VSS VDD  n8 n118 BUFx3_ASAP7_75t_L
XU72 VSS VDD  n118 result[6] INVx3_ASAP7_75t_L
XU73 VSS VDD  n120 result[2] INVx3_ASAP7_75t_L
XU74 VSS VDD  n119 result[4] INVx3_ASAP7_75t_L
XU75 VSS VDD  n10 n117 BUFx3_ASAP7_75t_L
XU76 VSS VDD  n117 result[8] INVx3_ASAP7_75t_L
XU77 VSS VDD  n12 n116 BUFx3_ASAP7_75t_L
XU78 VSS VDD  n116 result[10] INVx3_ASAP7_75t_L
XU79 VSS VDD  partial_sum[10] n106 INVx6_ASAP7_75t_L
XU80 VSS VDD  partial_sum[8] n95 INVx6_ASAP7_75t_L
XU81 VSS VDD  partial_sum[6] n84 INVx6_ASAP7_75t_L
XU82 VSS VDD  partial_sum[4] n73 INVx6_ASAP7_75t_L
XU83 VSS VDD  in_valid n51 INVx4_ASAP7_75t_L
XU84 VSS VDD  in_valid n52 INVx4_ASAP7_75t_L
XU85 VSS VDD  in_valid n115 INVx4_ASAP7_75t_L
XU86 VSS VDD  rst_n n53 INVx6_ASAP7_75t_L
XU87 VSS VDD  rst_n n54 INVx6_ASAP7_75t_L
XU88 VSS VDD  rst_n n55 INVx6_ASAP7_75t_L
XU89 VSS VDD  rst_n n56 INVx6_ASAP7_75t_L
XU90 VSS VDD  rst_n n15 INVx6_ASAP7_75t_L
XU91 VSS VDD  n2 TIELOx1_ASAP7_75t_L
XU92 VSS VDD  n14 result[12] INVxp33_ASAP7_75t_L
XU93 VSS VDD  n31 result[11] INVxp33_ASAP7_75t_L
XU94 VSS VDD  in_valid partial_sum[0] N_18 AND2x2_ASAP7_75t_L
XU95 VSS VDD  result[0] partial_sum[1] n57 NOR2xp33_ASAP7_75t_L
XU96 VSS VDD  n57 n48 n19 N_19 NOR3xp33_ASAP7_75t_L
XU97 VSS VDD  result[1] partial_sum[2] n59 NOR2xp33_ASAP7_75t_L
XU98 VSS VDD  n37 n34 n58 NOR2xp33_ASAP7_75t_L
XU99 VSS VDD  n59 n58 n60 NOR2xp33_ASAP7_75t_L
XU100 VSS VDD  n60 n48 A0  n61 HAxp5_ASAP7_75t_L
XU101 VSS VDD  n18 n61 N_20 NOR2xp33_ASAP7_75t_L
XU102 VSS VDD  n37 n62 n63 n68 MAJIxp5_ASAP7_75t_L
XU103 VSS VDD  result[2] partial_sum[3] n65 AND2x2_ASAP7_75t_L
XU104 VSS VDD  result[2] partial_sum[3] n64 NOR2xp33_ASAP7_75t_L
XU105 VSS VDD  n65 n64 n66 NOR2xp33_ASAP7_75t_L
XU106 VSS VDD  n68 n66 A1  n67 HAxp5_ASAP7_75t_L
XU107 VSS VDD  n21 n67 N_21 NOR2xp33_ASAP7_75t_L
XU108 VSS VDD  result[2] partial_sum[3] n68 n74 MAJIxp5_ASAP7_75t_L
XU109 VSS VDD  n38 n47 n70 NOR2xp33_ASAP7_75t_L
XU110 VSS VDD  result[3] partial_sum[4] n69 NOR2xp33_ASAP7_75t_L
XU111 VSS VDD  n70 n69 n71 NOR2xp33_ASAP7_75t_L
XU112 VSS VDD  n74 n71 n72 XOR2xp5_ASAP7_75t_L
XU113 VSS VDD  n51 n72 N_22 NOR2xp33_ASAP7_75t_L
XU114 VSS VDD  n38 n74 n73 n79 MAJIxp5_ASAP7_75t_L
XU115 VSS VDD  result[4] partial_sum[5] n76 AND2x2_ASAP7_75t_L
XU116 VSS VDD  result[4] partial_sum[5] n75 NOR2xp33_ASAP7_75t_L
XU117 VSS VDD  n76 n75 n77 NOR2xp33_ASAP7_75t_L
XU118 VSS VDD  n79 n77 A2  n78 HAxp5_ASAP7_75t_L
XU119 VSS VDD  n49 n78 N_23 NOR2xp33_ASAP7_75t_L
XU120 VSS VDD  result[4] partial_sum[5] n79 n85 MAJIxp5_ASAP7_75t_L
XU121 VSS VDD  n39 n46 n81 NOR2xp33_ASAP7_75t_L
XU122 VSS VDD  result[5] partial_sum[6] n80 NOR2xp33_ASAP7_75t_L
XU123 VSS VDD  n81 n80 n82 NOR2xp33_ASAP7_75t_L
XU124 VSS VDD  n85 n82 n83 XOR2xp5_ASAP7_75t_L
XU125 VSS VDD  n16 n83 N_24 NOR2xp33_ASAP7_75t_L
XU126 VSS VDD  n39 n85 n84 n90 MAJIxp5_ASAP7_75t_L
XU127 VSS VDD  result[6] partial_sum[7] n87 AND2x2_ASAP7_75t_L
XU128 VSS VDD  result[6] partial_sum[7] n86 NOR2xp33_ASAP7_75t_L
XU129 VSS VDD  n87 n86 n88 NOR2xp33_ASAP7_75t_L
XU130 VSS VDD  n90 n88 A3  n89 HAxp5_ASAP7_75t_L
XU131 VSS VDD  n52 n89 N_25 NOR2xp33_ASAP7_75t_L
XU132 VSS VDD  result[6] partial_sum[7] n90 n96 MAJIxp5_ASAP7_75t_L
XU133 VSS VDD  n32 n45 n92 NOR2xp33_ASAP7_75t_L
XU134 VSS VDD  result[7] partial_sum[8] n91 NOR2xp33_ASAP7_75t_L
XU135 VSS VDD  n92 n91 n93 NOR2xp33_ASAP7_75t_L
XU136 VSS VDD  n96 n93 n94 XOR2xp5_ASAP7_75t_L
XU137 VSS VDD  n115 n94 N_26 NOR2xp33_ASAP7_75t_L
XU138 VSS VDD  n32 n96 n95 n101 MAJIxp5_ASAP7_75t_L
XU139 VSS VDD  result[8] partial_sum[9] n98 AND2x2_ASAP7_75t_L
XU140 VSS VDD  result[8] partial_sum[9] n97 NOR2xp33_ASAP7_75t_L
XU141 VSS VDD  n98 n97 n99 NOR2xp33_ASAP7_75t_L
XU142 VSS VDD  n101 n99 A4  n100 HAxp5_ASAP7_75t_L
XU143 VSS VDD  n50 n100 N_27 NOR2xp33_ASAP7_75t_L
XU144 VSS VDD  result[8] partial_sum[9] n101 n107 MAJIxp5_ASAP7_75t_L
XU145 VSS VDD  n33 n44 n103 NOR2xp33_ASAP7_75t_L
XU146 VSS VDD  result[9] partial_sum[10] n102 NOR2xp33_ASAP7_75t_L
XU147 VSS VDD  n103 n102 n104 NOR2xp33_ASAP7_75t_L
XU148 VSS VDD  n107 n104 n105 XOR2xp5_ASAP7_75t_L
XU149 VSS VDD  n17 n105 N_28 NOR2xp33_ASAP7_75t_L
XU150 VSS VDD  n33 n107 n106 n112 MAJIxp5_ASAP7_75t_L
XU151 VSS VDD  result[10] partial_sum[11] n109 NOR2xp33_ASAP7_75t_L
XU152 VSS VDD  result[10] partial_sum[11] n108 AND2x2_ASAP7_75t_L
XU153 VSS VDD  n109 n108 n110 NOR2xp33_ASAP7_75t_L
XU154 VSS VDD  n112 n110 A5  n111 HAxp5_ASAP7_75t_L
XU155 VSS VDD  n22 n111 N_29 NOR2xp33_ASAP7_75t_L
XU156 VSS VDD  result[10] partial_sum[11] n112 n113 MAJIxp5_ASAP7_75t_L
XU157 VSS VDD  partial_sum[12] n113 n31 A6  n114 FAx1_ASAP7_75t_L
XU158 VSS VDD  n20 n114 N_30 NOR2xp33_ASAP7_75t_L
.ENDS


