.TITLE DIC_Final

***-----------------------***
***        setting        ***
***-----------------------***

.protect
.include '../08_TECH/LIB/7nm_TT.pm'
.include '../08_TECH/LIB/16mos.pm'
.include '../08_TECH/LIB/asap7sc7p5t_SIMPLE_RVT.sp' 
.include '../08_TECH/LIB/asap7sc7p5t_SEQ_RVT.sp'    
.include '../08_TECH/LIB/asap7sc7p5t_INVBUF_RVT.sp' 
.include '../08_TECH/LIB/asap7sc7p5t_AO_RVT.sp'     
.include '../08_TECH/LIB/asap7sc7p5t_OA_RVT.sp'     
.include './Adder_tree_SYN_new.sp'
.include './Accumulator_SYN_new.sp'
.unprotect

.VEC "mul.vec" 

*** Voltage: 0.7V ***
.PARAM supply=0.7v

*** Temperature: 25C ***
.TEMP 25

***********************************
* Transition Analysis             *
***********************************
.TRAN 1ps 20ns 

***********************************
* HSPICE Options                  *
***********************************
.OPTION POST PROBE
.OPTION NOMOD BRIEF MEASDGT=7 
.OPTION CAPTAB NOTOP AUTOSTOP

***********************************
* Output Signals                  *
***********************************
.probe tran v(*) i(*)


***********************************
* Define Global Nets              *
***********************************
.GLOBAL VDD GND BL BLB

***********************************
* Voltage Sources                 *
***********************************
vdd     VDD   0  DC supply
vss     VSS   0  DC 0
vbl     BL    0   DC supply/2
vblb    BLB   0   DC supply/2

***********************************
* Measurement Commands            *
***********************************
.meas pwr avg POWER



***-----------------------***
***        circuit        ***
***-----------------------***


* // Xbuf Input In_bar INV
* // ADD INPUT BUFFER
* // WEIGHT IS INITIALIZE IN THE SRAM
* // SO CIM OPERATION IS READ THE WEIGHT AND THEN DO DOT PRODUCT 
* XI11 I111 I111_inv INV
* XI12 I112 I112_inv INV
* XI13 I113 I113_inv INV
* XI14 I114 I114_inv INV
* XI15 I121 I121_inv INV
* XI16 I122 I122_inv INV
* XI17 I123 I123_inv INV
* XI18 I124 I124_inv INV
* XI19 I131 I131_inv INV
* XI20 I132 I132_inv INV
* XI21 I133 I133_inv INV
* XI22 I134 I134_inv INV
* XI23 I141 I141_inv INV
* XI24 I142 I142_inv INV
* XI25 I143 I143_inv INV
* XI26 I144 I144_inv INV
* XI27 I151 I151_inv INV
* XI28 I152 I152_inv INV
* XI29 I153 I153_inv INV
* XI30 I154 I154_inv INV
* XI31 I161 I161_inv INV
* XI32 I162 I162_inv INV
* XI33 I163 I163_inv INV
* XI34 I164 I164_inv INV
* XI35 I171 I171_inv INV
* XI36 I172 I172_inv INV
* XI37 I173 I173_inv INV
* XI38 I174 I174_inv INV
* XI39 I181 I181_inv INV
* XI40 I182 I182_inv INV
* XI41 I183 I183_inv INV
* XI42 I184 I184_inv INV
* XI43 I191 I191_inv INV
* XI44 I192 I192_inv INV
* XI45 I193 I193_inv INV
* XI46 I194 I194_inv INV
* XI47 I1101 I1101_inv INV
* XI48 I1102 I1102_inv INV
* XI49 I1103 I1103_inv INV
* XI50 I1104 I1104_inv INV
* XI51 I1111 I1111_inv INV
* XI52 I1112 I1112_inv INV
* XI53 I1113 I1113_inv INV
* XI54 I1114 I1114_inv INV
* XI55 I1121 I1121_inv INV
* XI56 I1122 I1122_inv INV
* XI57 I1123 I1123_inv INV
* XI58 I1124 I1124_inv INV
* XI59 I1131 I1131_inv INV
* XI60 I1132 I1132_inv INV
* XI61 I1133 I1133_inv INV
* XI62 I1134 I1134_inv INV
* XI63 I1141 I1141_inv INV
* XI64 I1142 I1142_inv INV
* XI65 I1143 I1143_inv INV
* XI66 I1144 I1144_inv INV
* XI67 I1151 I1151_inv INV
* XI68 I1152 I1152_inv INV
* XI69 I1153 I1153_inv INV
* XI70 I1154 I1154_inv INV
* XI71 I1161 I1161_inv INV
* XI72 I1162 I1162_inv INV
* XI73 I1163 I1163_inv INV
* XI74 I1164 I1164_inv INV
* XI75 I1171 I1171_inv INV
* XI76 I1172 I1172_inv INV
* XI77 I1173 I1173_inv INV
* XI78 I1174 I1174_inv INV
* XI79 I1181 I1181_inv INV
* XI80 I1182 I1182_inv INV
* XI81 I1183 I1183_inv INV
* XI82 I1184 I1184_inv INV
* XI83 I1191 I1191_inv INV
* XI84 I1192 I1192_inv INV
* XI85 I1193 I1193_inv INV
* XI86 I1194 I1194_inv INV
* XI87 I1201 I1201_inv INV
* XI88 I1202 I1202_inv INV
* XI89 I1203 I1203_inv INV
* XI90 I1204 I1204_inv INV
* XI91 I1211 I1211_inv INV
* XI92 I1212 I1212_inv INV
* XI93 I1213 I1213_inv INV
* XI94 I1214 I1214_inv INV
* XI95 I1221 I1221_inv INV
* XI96 I1222 I1222_inv INV
* XI97 I1223 I1223_inv INV
* XI98 I1224 I1224_inv INV
* XI99 I1231 I1231_inv INV
* XI100 I1232 I1232_inv INV
* XI101 I1233 I1233_inv INV
* XI102 I1234 I1234_inv INV
* XI103 I1241 I1241_inv INV
* XI104 I1242 I1242_inv INV
* XI105 I1243 I1243_inv INV
* XI106 I1244 I1244_inv INV
* XI107 I1251 I1251_inv INV
* XI108 I1252 I1252_inv INV
* XI109 I1253 I1253_inv INV
* XI110 I1254 I1254_inv INV
* XI111 I1261 I1261_inv INV
* XI112 I1262 I1262_inv INV
* XI113 I1263 I1263_inv INV
* XI114 I1264 I1264_inv INV
* XI115 I1271 I1271_inv INV
* XI116 I1272 I1272_inv INV
* XI117 I1273 I1273_inv INV
* XI118 I1274 I1274_inv INV
* XI119 I1281 I1281_inv INV
* XI120 I1282 I1282_inv INV
* XI121 I1283 I1283_inv INV
* XI122 I1284 I1284_inv INV
* XI123 I1291 I1291_inv INV
* XI124 I1292 I1292_inv INV
* XI125 I1293 I1293_inv INV
* XI126 I1294 I1294_inv INV
* XI127 I1301 I1301_inv INV
* XI128 I1302 I1302_inv INV
* XI129 I1303 I1303_inv INV
* XI130 I1304 I1304_inv INV
* XI131 I1311 I1311_inv INV
* XI132 I1312 I1312_inv INV
* XI133 I1313 I1313_inv INV
* XI134 I1314 I1314_inv INV
* XI135 I1321 I1321_inv INV
* XI136 I1322 I1322_inv INV
* XI137 I1323 I1323_inv INV
* XI138 I1324 I1324_inv INV
* XI139 I211 I211_inv INV
* XI140 I212 I212_inv INV
* XI141 I213 I213_inv INV
* XI142 I214 I214_inv INV
* XI143 I221 I221_inv INV
* XI144 I222 I222_inv INV
* XI145 I223 I223_inv INV
* XI146 I224 I224_inv INV
* XI147 I231 I231_inv INV
* XI148 I232 I232_inv INV
* XI149 I233 I233_inv INV
* XI150 I234 I234_inv INV
* XI151 I241 I241_inv INV
* XI152 I242 I242_inv INV
* XI153 I243 I243_inv INV
* XI154 I244 I244_inv INV
* XI155 I251 I251_inv INV
* XI156 I252 I252_inv INV
* XI157 I253 I253_inv INV
* XI158 I254 I254_inv INV
* XI159 I261 I261_inv INV
* XI160 I262 I262_inv INV
* XI161 I263 I263_inv INV
* XI162 I264 I264_inv INV
* XI163 I271 I271_inv INV
* XI164 I272 I272_inv INV
* XI165 I273 I273_inv INV
* XI166 I274 I274_inv INV
* XI167 I281 I281_inv INV
* XI168 I282 I282_inv INV
* XI169 I283 I283_inv INV
* XI170 I284 I284_inv INV
* XI171 I291 I291_inv INV
* XI172 I292 I292_inv INV
* XI173 I293 I293_inv INV
* XI174 I294 I294_inv INV
* XI175 I2101 I2101_inv INV
* XI176 I2102 I2102_inv INV
* XI177 I2103 I2103_inv INV
* XI178 I2104 I2104_inv INV
* XI179 I2111 I2111_inv INV
* XI180 I2112 I2112_inv INV
* XI181 I2113 I2113_inv INV
* XI182 I2114 I2114_inv INV
* XI183 I2121 I2121_inv INV
* XI184 I2122 I2122_inv INV
* XI185 I2123 I2123_inv INV
* XI186 I2124 I2124_inv INV
* XI187 I2131 I2131_inv INV
* XI188 I2132 I2132_inv INV
* XI189 I2133 I2133_inv INV
* XI190 I2134 I2134_inv INV
* XI191 I2141 I2141_inv INV
* XI192 I2142 I2142_inv INV
* XI193 I2143 I2143_inv INV
* XI194 I2144 I2144_inv INV
* XI195 I2151 I2151_inv INV
* XI196 I2152 I2152_inv INV
* XI197 I2153 I2153_inv INV
* XI198 I2154 I2154_inv INV
* XI199 I2161 I2161_inv INV
* XI200 I2162 I2162_inv INV
* XI201 I2163 I2163_inv INV
* XI202 I2164 I2164_inv INV
* XI203 I2171 I2171_inv INV
* XI204 I2172 I2172_inv INV
* XI205 I2173 I2173_inv INV
* XI206 I2174 I2174_inv INV
* XI207 I2181 I2181_inv INV
* XI208 I2182 I2182_inv INV
* XI209 I2183 I2183_inv INV
* XI210 I2184 I2184_inv INV
* XI211 I2191 I2191_inv INV
* XI212 I2192 I2192_inv INV
* XI213 I2193 I2193_inv INV
* XI214 I2194 I2194_inv INV
* XI215 I2201 I2201_inv INV
* XI216 I2202 I2202_inv INV
* XI217 I2203 I2203_inv INV
* XI218 I2204 I2204_inv INV
* XI219 I2211 I2211_inv INV
* XI220 I2212 I2212_inv INV
* XI221 I2213 I2213_inv INV
* XI222 I2214 I2214_inv INV
* XI223 I2221 I2221_inv INV
* XI224 I2222 I2222_inv INV
* XI225 I2223 I2223_inv INV
* XI226 I2224 I2224_inv INV
* XI227 I2231 I2231_inv INV
* XI228 I2232 I2232_inv INV
* XI229 I2233 I2233_inv INV
* XI230 I2234 I2234_inv INV
* XI231 I2241 I2241_inv INV
* XI232 I2242 I2242_inv INV
* XI233 I2243 I2243_inv INV
* XI234 I2244 I2244_inv INV
* XI235 I2251 I2251_inv INV
* XI236 I2252 I2252_inv INV
* XI237 I2253 I2253_inv INV
* XI238 I2254 I2254_inv INV
* XI239 I2261 I2261_inv INV
* XI240 I2262 I2262_inv INV
* XI241 I2263 I2263_inv INV
* XI242 I2264 I2264_inv INV
* XI243 I2271 I2271_inv INV
* XI244 I2272 I2272_inv INV
* XI245 I2273 I2273_inv INV
* XI246 I2274 I2274_inv INV
* XI247 I2281 I2281_inv INV
* XI248 I2282 I2282_inv INV
* XI249 I2283 I2283_inv INV
* XI250 I2284 I2284_inv INV
* XI251 I2291 I2291_inv INV
* XI252 I2292 I2292_inv INV
* XI253 I2293 I2293_inv INV
* XI254 I2294 I2294_inv INV
* XI255 I2301 I2301_inv INV
* XI256 I2302 I2302_inv INV
* XI257 I2303 I2303_inv INV
* XI258 I2304 I2304_inv INV
* XI259 I2311 I2311_inv INV
* XI260 I2312 I2312_inv INV
* XI261 I2313 I2313_inv INV
* XI262 I2314 I2314_inv INV
* XI263 I2321 I2321_inv INV
* XI264 I2322 I2322_inv INV
* XI265 I2323 I2323_inv INV
* XI266 I2324 I2324_inv INV
* XI267 I311 I311_inv INV
* XI268 I312 I312_inv INV
* XI269 I313 I313_inv INV
* XI270 I314 I314_inv INV
* XI271 I321 I321_inv INV
* XI272 I322 I322_inv INV
* XI273 I323 I323_inv INV
* XI274 I324 I324_inv INV
* XI275 I331 I331_inv INV
* XI276 I332 I332_inv INV
* XI277 I333 I333_inv INV
* XI278 I334 I334_inv INV
* XI279 I341 I341_inv INV
* XI280 I342 I342_inv INV
* XI281 I343 I343_inv INV
* XI282 I344 I344_inv INV
* XI283 I351 I351_inv INV
* XI284 I352 I352_inv INV
* XI285 I353 I353_inv INV
* XI286 I354 I354_inv INV
* XI287 I361 I361_inv INV
* XI288 I362 I362_inv INV
* XI289 I363 I363_inv INV
* XI290 I364 I364_inv INV
* XI291 I371 I371_inv INV
* XI292 I372 I372_inv INV
* XI293 I373 I373_inv INV
* XI294 I374 I374_inv INV
* XI295 I381 I381_inv INV
* XI296 I382 I382_inv INV
* XI297 I383 I383_inv INV
* XI298 I384 I384_inv INV
* XI299 I391 I391_inv INV
* XI300 I392 I392_inv INV
* XI301 I393 I393_inv INV
* XI302 I394 I394_inv INV
* XI303 I3101 I3101_inv INV
* XI304 I3102 I3102_inv INV
* XI305 I3103 I3103_inv INV
* XI306 I3104 I3104_inv INV
* XI307 I3111 I3111_inv INV
* XI308 I3112 I3112_inv INV
* XI309 I3113 I3113_inv INV
* XI310 I3114 I3114_inv INV
* XI311 I3121 I3121_inv INV
* XI312 I3122 I3122_inv INV
* XI313 I3123 I3123_inv INV
* XI314 I3124 I3124_inv INV
* XI315 I3131 I3131_inv INV
* XI316 I3132 I3132_inv INV
* XI317 I3133 I3133_inv INV
* XI318 I3134 I3134_inv INV
* XI319 I3141 I3141_inv INV
* XI320 I3142 I3142_inv INV
* XI321 I3143 I3143_inv INV
* XI322 I3144 I3144_inv INV
* XI323 I3151 I3151_inv INV
* XI324 I3152 I3152_inv INV
* XI325 I3153 I3153_inv INV
* XI326 I3154 I3154_inv INV
* XI327 I3161 I3161_inv INV
* XI328 I3162 I3162_inv INV
* XI329 I3163 I3163_inv INV
* XI330 I3164 I3164_inv INV
* XI331 I3171 I3171_inv INV
* XI332 I3172 I3172_inv INV
* XI333 I3173 I3173_inv INV
* XI334 I3174 I3174_inv INV
* XI335 I3181 I3181_inv INV
* XI336 I3182 I3182_inv INV
* XI337 I3183 I3183_inv INV
* XI338 I3184 I3184_inv INV
* XI339 I3191 I3191_inv INV
* XI340 I3192 I3192_inv INV
* XI341 I3193 I3193_inv INV
* XI342 I3194 I3194_inv INV
* XI343 I3201 I3201_inv INV
* XI344 I3202 I3202_inv INV
* XI345 I3203 I3203_inv INV
* XI346 I3204 I3204_inv INV
* XI347 I3211 I3211_inv INV
* XI348 I3212 I3212_inv INV
* XI349 I3213 I3213_inv INV
* XI350 I3214 I3214_inv INV
* XI351 I3221 I3221_inv INV
* XI352 I3222 I3222_inv INV
* XI353 I3223 I3223_inv INV
* XI354 I3224 I3224_inv INV
* XI355 I3231 I3231_inv INV
* XI356 I3232 I3232_inv INV
* XI357 I3233 I3233_inv INV
* XI358 I3234 I3234_inv INV
* XI359 I3241 I3241_inv INV
* XI360 I3242 I3242_inv INV
* XI361 I3243 I3243_inv INV
* XI362 I3244 I3244_inv INV
* XI363 I3251 I3251_inv INV
* XI364 I3252 I3252_inv INV
* XI365 I3253 I3253_inv INV
* XI366 I3254 I3254_inv INV
* XI367 I3261 I3261_inv INV
* XI368 I3262 I3262_inv INV
* XI369 I3263 I3263_inv INV
* XI370 I3264 I3264_inv INV
* XI371 I3271 I3271_inv INV
* XI372 I3272 I3272_inv INV
* XI373 I3273 I3273_inv INV
* XI374 I3274 I3274_inv INV
* XI375 I3281 I3281_inv INV
* XI376 I3282 I3282_inv INV
* XI377 I3283 I3283_inv INV
* XI378 I3284 I3284_inv INV
* XI379 I3291 I3291_inv INV
* XI380 I3292 I3292_inv INV
* XI381 I3293 I3293_inv INV
* XI382 I3294 I3294_inv INV
* XI383 I3301 I3301_inv INV
* XI384 I3302 I3302_inv INV
* XI385 I3303 I3303_inv INV
* XI386 I3304 I3304_inv INV
* XI387 I3311 I3311_inv INV
* XI388 I3312 I3312_inv INV
* XI389 I3313 I3313_inv INV
* XI390 I3314 I3314_inv INV
* XI391 I3321 I3321_inv INV
* XI392 I3322 I3322_inv INV
* XI393 I3323 I3323_inv INV
* XI394 I3324 I3324_inv INV
* XI395 I411 I411_inv INV
* XI396 I412 I412_inv INV
* XI397 I413 I413_inv INV
* XI398 I414 I414_inv INV
* XI399 I421 I421_inv INV
* XI400 I422 I422_inv INV
* XI401 I423 I423_inv INV
* XI402 I424 I424_inv INV
* XI403 I431 I431_inv INV
* XI404 I432 I432_inv INV
* XI405 I433 I433_inv INV
* XI406 I434 I434_inv INV
* XI407 I441 I441_inv INV
* XI408 I442 I442_inv INV
* XI409 I443 I443_inv INV
* XI410 I444 I444_inv INV
* XI411 I451 I451_inv INV
* XI412 I452 I452_inv INV
* XI413 I453 I453_inv INV
* XI414 I454 I454_inv INV
* XI415 I461 I461_inv INV
* XI416 I462 I462_inv INV
* XI417 I463 I463_inv INV
* XI418 I464 I464_inv INV
* XI419 I471 I471_inv INV
* XI420 I472 I472_inv INV
* XI421 I473 I473_inv INV
* XI422 I474 I474_inv INV
* XI423 I481 I481_inv INV
* XI424 I482 I482_inv INV
* XI425 I483 I483_inv INV
* XI426 I484 I484_inv INV
* XI427 I491 I491_inv INV
* XI428 I492 I492_inv INV
* XI429 I493 I493_inv INV
* XI430 I494 I494_inv INV
* XI431 I4101 I4101_inv INV
* XI432 I4102 I4102_inv INV
* XI433 I4103 I4103_inv INV
* XI434 I4104 I4104_inv INV
* XI435 I4111 I4111_inv INV
* XI436 I4112 I4112_inv INV
* XI437 I4113 I4113_inv INV
* XI438 I4114 I4114_inv INV
* XI439 I4121 I4121_inv INV
* XI440 I4122 I4122_inv INV
* XI441 I4123 I4123_inv INV
* XI442 I4124 I4124_inv INV
* XI443 I4131 I4131_inv INV
* XI444 I4132 I4132_inv INV
* XI445 I4133 I4133_inv INV
* XI446 I4134 I4134_inv INV
* XI447 I4141 I4141_inv INV
* XI448 I4142 I4142_inv INV
* XI449 I4143 I4143_inv INV
* XI450 I4144 I4144_inv INV
* XI451 I4151 I4151_inv INV
* XI452 I4152 I4152_inv INV
* XI453 I4153 I4153_inv INV
* XI454 I4154 I4154_inv INV
* XI455 I4161 I4161_inv INV
* XI456 I4162 I4162_inv INV
* XI457 I4163 I4163_inv INV
* XI458 I4164 I4164_inv INV
* XI459 I4171 I4171_inv INV
* XI460 I4172 I4172_inv INV
* XI461 I4173 I4173_inv INV
* XI462 I4174 I4174_inv INV
* XI463 I4181 I4181_inv INV
* XI464 I4182 I4182_inv INV
* XI465 I4183 I4183_inv INV
* XI466 I4184 I4184_inv INV
* XI467 I4191 I4191_inv INV
* XI468 I4192 I4192_inv INV
* XI469 I4193 I4193_inv INV
* XI470 I4194 I4194_inv INV
* XI471 I4201 I4201_inv INV
* XI472 I4202 I4202_inv INV
* XI473 I4203 I4203_inv INV
* XI474 I4204 I4204_inv INV
* XI475 I4211 I4211_inv INV
* XI476 I4212 I4212_inv INV
* XI477 I4213 I4213_inv INV
* XI478 I4214 I4214_inv INV
* XI479 I4221 I4221_inv INV
* XI480 I4222 I4222_inv INV
* XI481 I4223 I4223_inv INV
* XI482 I4224 I4224_inv INV
* XI483 I4231 I4231_inv INV
* XI484 I4232 I4232_inv INV
* XI485 I4233 I4233_inv INV
* XI486 I4234 I4234_inv INV
* XI487 I4241 I4241_inv INV
* XI488 I4242 I4242_inv INV
* XI489 I4243 I4243_inv INV
* XI490 I4244 I4244_inv INV
* XI491 I4251 I4251_inv INV
* XI492 I4252 I4252_inv INV
* XI493 I4253 I4253_inv INV
* XI494 I4254 I4254_inv INV
* XI495 I4261 I4261_inv INV
* XI496 I4262 I4262_inv INV
* XI497 I4263 I4263_inv INV
* XI498 I4264 I4264_inv INV
* XI499 I4271 I4271_inv INV
* XI500 I4272 I4272_inv INV
* XI501 I4273 I4273_inv INV
* XI502 I4274 I4274_inv INV
* XI503 I4281 I4281_inv INV
* XI504 I4282 I4282_inv INV
* XI505 I4283 I4283_inv INV
* XI506 I4284 I4284_inv INV
* XI507 I4291 I4291_inv INV
* XI508 I4292 I4292_inv INV
* XI509 I4293 I4293_inv INV
* XI510 I4294 I4294_inv INV
* XI511 I4301 I4301_inv INV
* XI512 I4302 I4302_inv INV
* XI513 I4303 I4303_inv INV
* XI514 I4304 I4304_inv INV
* XI515 I4311 I4311_inv INV
* XI516 I4312 I4312_inv INV
* XI517 I4313 I4313_inv INV
* XI518 I4314 I4314_inv INV
* XI519 I4321 I4321_inv INV
* XI520 I4322 I4322_inv INV
* XI521 I4323 I4323_inv INV
* XI522 I4324 I4324_inv INV

XI11 I11 I11_buf INV
XB11 I11_buf I11_inv Buffer

XI15 I12 I12_buf INV
XB15 I12_buf I12_inv Buffer

XI19 I13 I13_buf INV
XB19 I13_buf I13_inv Buffer

XI23 I14 I14_buf INV
XB23 I14_buf I14_inv Buffer

XI27 I15 I15_buf INV
XB27 I15_buf I15_inv Buffer

XI31 I16 I16_buf INV
XB31 I16_buf I16_inv Buffer

XI35 I17 I17_buf INV
XB35 I17_buf I17_inv Buffer

XI39 I18 I18_buf INV
XB39 I18_buf I18_inv Buffer

XI43 I19 I19_buf INV
XB43 I19_buf I19_inv Buffer

XI47 I110 I110_buf INV
XB47 I110_buf I110_inv Buffer

XI51 I111 I111_buf INV
XB51 I111_buf I111_inv Buffer

XI55 I112 I112_buf INV
XB55 I112_buf I112_inv Buffer

XI59 I113 I113_buf INV
XB59 I113_buf I113_inv Buffer

XI63 I114 I114_buf INV
XB63 I114_buf I114_inv Buffer

XI67 I115 I115_buf INV
XB67 I115_buf I115_inv Buffer

XI71 I116 I116_buf INV
XB71 I116_buf I116_inv Buffer

XI75 I117 I117_buf INV
XB75 I117_buf I117_inv Buffer

XI79 I118 I118_buf INV
XB79 I118_buf I118_inv Buffer

XI83 I119 I119_buf INV
XB83 I119_buf I119_inv Buffer

XI87 I120 I120_buf INV
XB87 I120_buf I120_inv Buffer

XI91 I121 I121_buf INV
XB91 I121_buf I121_inv Buffer

XI95 I122 I122_buf INV
XB95 I122_buf I122_inv Buffer

XI99 I123 I123_buf INV
XB99 I123_buf I123_inv Buffer

XI103 I124 I124_buf INV
XB103 I124_buf I124_inv Buffer

XI107 I125 I125_buf INV
XB107 I125_buf I125_inv Buffer

XI111 I126 I126_buf INV
XB111 I126_buf I126_inv Buffer

XI115 I127 I127_buf INV
XB115 I127_buf I127_inv Buffer

XI119 I128 I128_buf INV
XB119 I128_buf I128_inv Buffer

XI123 I129 I129_buf INV
XB123 I129_buf I129_inv Buffer

XI127 I130 I130_buf INV
XB127 I130_buf I130_inv Buffer

XI131 I131 I131_buf INV
XB131 I131_buf I131_inv Buffer

XI135 I132 I132_buf INV
XB135 I132_buf I132_inv Buffer

XI139 I21 I21_buf INV
XB139 I21_buf I21_inv Buffer

XI143 I22 I22_buf INV
XB143 I22_buf I22_inv Buffer

XI147 I23 I23_buf INV
XB147 I23_buf I23_inv Buffer

XI151 I24 I24_buf INV
XB151 I24_buf I24_inv Buffer

XI155 I25 I25_buf INV
XB155 I25_buf I25_inv Buffer

XI159 I26 I26_buf INV
XB159 I26_buf I26_inv Buffer

XI163 I27 I27_buf INV
XB163 I27_buf I27_inv Buffer

XI167 I28 I28_buf INV
XB167 I28_buf I28_inv Buffer

XI171 I29 I29_buf INV
XB171 I29_buf I29_inv Buffer

XI175 I210 I210_buf INV
XB175 I210_buf I210_inv Buffer

XI179 I211 I211_buf INV
XB179 I211_buf I211_inv Buffer

XI183 I212 I212_buf INV
XB183 I212_buf I212_inv Buffer

XI187 I213 I213_buf INV
XB187 I213_buf I213_inv Buffer

XI191 I214 I214_buf INV
XB191 I214_buf I214_inv Buffer

XI195 I215 I215_buf INV
XB195 I215_buf I215_inv Buffer

XI199 I216 I216_buf INV
XB199 I216_buf I216_inv Buffer

XI203 I217 I217_buf INV
XB203 I217_buf I217_inv Buffer

XI207 I218 I218_buf INV
XB207 I218_buf I218_inv Buffer

XI211 I219 I219_buf INV
XB211 I219_buf I219_inv Buffer

XI215 I220 I220_buf INV
XB215 I220_buf I220_inv Buffer

XI219 I221 I221_buf INV
XB219 I221_buf I221_inv Buffer

XI223 I222 I222_buf INV
XB223 I222_buf I222_inv Buffer

XI227 I223 I223_buf INV
XB227 I223_buf I223_inv Buffer

XI231 I224 I224_buf INV
XB231 I224_buf I224_inv Buffer

XI235 I225 I225_buf INV
XB235 I225_buf I225_inv Buffer

XI239 I226 I226_buf INV
XB239 I226_buf I226_inv Buffer

XI243 I227 I227_buf INV
XB243 I227_buf I227_inv Buffer

XI247 I228 I228_buf INV
XB247 I228_buf I228_inv Buffer

XI251 I229 I229_buf INV
XB251 I229_buf I229_inv Buffer

XI255 I230 I230_buf INV
XB255 I230_buf I230_inv Buffer

XI259 I231 I231_buf INV
XB259 I231_buf I231_inv Buffer

XI263 I232 I232_buf INV
XB263 I232_buf I232_inv Buffer

XI267 I31 I31_buf INV
XB267 I31_buf I31_inv Buffer

XI271 I32 I32_buf INV
XB271 I32_buf I32_inv Buffer

XI275 I33 I33_buf INV
XB275 I33_buf I33_inv Buffer

XI279 I34 I34_buf INV
XB279 I34_buf I34_inv Buffer

XI283 I35 I35_buf INV
XB283 I35_buf I35_inv Buffer

XI287 I36 I36_buf INV
XB287 I36_buf I36_inv Buffer

XI291 I37 I37_buf INV
XB291 I37_buf I37_inv Buffer

XI295 I38 I38_buf INV
XB295 I38_buf I38_inv Buffer

XI299 I39 I39_buf INV
XB299 I39_buf I39_inv Buffer

XI303 I310 I310_buf INV
XB303 I310_buf I310_inv Buffer

XI307 I311 I311_buf INV
XB307 I311_buf I311_inv Buffer

XI311 I312 I312_buf INV
XB311 I312_buf I312_inv Buffer

XI315 I313 I313_buf INV
XB315 I313_buf I313_inv Buffer

XI319 I314 I314_buf INV
XB319 I314_buf I314_inv Buffer

XI323 I315 I315_buf INV
XB323 I315_buf I315_inv Buffer

XI327 I316 I316_buf INV
XB327 I316_buf I316_inv Buffer

XI331 I317 I317_buf INV
XB331 I317_buf I317_inv Buffer

XI335 I318 I318_buf INV
XB335 I318_buf I318_inv Buffer

XI339 I319 I319_buf INV
XB339 I319_buf I319_inv Buffer

XI343 I320 I320_buf INV
XB343 I320_buf I320_inv Buffer

XI347 I321 I321_buf INV
XB347 I321_buf I321_inv Buffer

XI351 I322 I322_buf INV
XB351 I322_buf I322_inv Buffer

XI355 I323 I323_buf INV
XB355 I323_buf I323_inv Buffer

XI359 I324 I324_buf INV
XB359 I324_buf I324_inv Buffer

XI363 I325 I325_buf INV
XB363 I325_buf I325_inv Buffer

XI367 I326 I326_buf INV
XB367 I326_buf I326_inv Buffer

XI371 I327 I327_buf INV
XB371 I327_buf I327_inv Buffer

XI375 I328 I328_buf INV
XB375 I328_buf I328_inv Buffer

XI379 I329 I329_buf INV
XB379 I329_buf I329_inv Buffer

XI383 I330 I330_buf INV
XB383 I330_buf I330_inv Buffer

XI387 I331 I331_buf INV
XB387 I331_buf I331_inv Buffer

XI391 I332 I332_buf INV
XB391 I332_buf I332_inv Buffer

XI395 I41 I41_buf INV
XB395 I41_buf I41_inv Buffer

XI399 I42 I42_buf INV
XB399 I42_buf I42_inv Buffer

XI403 I43 I43_buf INV
XB403 I43_buf I43_inv Buffer

XI407 I44 I44_buf INV
XB407 I44_buf I44_inv Buffer

XI411 I45 I45_buf INV
XB411 I45_buf I45_inv Buffer

XI415 I46 I46_buf INV
XB415 I46_buf I46_inv Buffer

XI419 I47 I47_buf INV
XB419 I47_buf I47_inv Buffer

XI423 I48 I48_buf INV
XB423 I48_buf I48_inv Buffer

XI427 I49 I49_buf INV
XB427 I49_buf I49_inv Buffer

XI431 I410 I410_buf INV
XB431 I410_buf I410_inv Buffer

XI435 I411 I411_buf INV
XB435 I411_buf I411_inv Buffer

XI439 I412 I412_buf INV
XB439 I412_buf I412_inv Buffer

XI443 I413 I413_buf INV
XB443 I413_buf I413_inv Buffer

XI447 I414 I414_buf INV
XB447 I414_buf I414_inv Buffer

XI451 I415 I415_buf INV
XB451 I415_buf I415_inv Buffer

XI455 I416 I416_buf INV
XB455 I416_buf I416_inv Buffer

XI459 I417 I417_buf INV
XB459 I417_buf I417_inv Buffer

XI463 I418 I418_buf INV
XB463 I418_buf I418_inv Buffer

XI467 I419 I419_buf INV
XB467 I419_buf I419_inv Buffer

XI471 I420 I420_buf INV
XB471 I420_buf I420_inv Buffer

XI475 I421 I421_buf INV
XB475 I421_buf I421_inv Buffer

XI479 I422 I422_buf INV
XB479 I422_buf I422_inv Buffer

XI483 I423 I423_buf INV
XB483 I423_buf I423_inv Buffer

XI487 I424 I424_buf INV
XB487 I424_buf I424_inv Buffer

XI491 I425 I425_buf INV
XB491 I425_buf I425_inv Buffer

XI495 I426 I426_buf INV
XB495 I426_buf I426_inv Buffer

XI499 I427 I427_buf INV
XB499 I427_buf I427_inv Buffer

XI503 I428 I428_buf INV
XB503 I428_buf I428_inv Buffer

XI507 I429 I429_buf INV
XB507 I429_buf I429_inv Buffer

XI511 I430 I430_buf INV
XB511 I430_buf I430_inv Buffer

XI515 I431 I431_buf INV
XB515 I431_buf I431_inv Buffer

XI519 I432 I432_buf INV
XB519 I432_buf I432_inv Buffer


X1 I11_inv O_1_1_1 WL_1_1 BL BLB W_1_1_1 W_1_1_1_bar CIM_cell
X2 I11_inv O_1_1_2 WL_1_2 BL BLB W_1_1_2 W_1_1_2_bar CIM_cell
X3 I11_inv O_1_1_3 WL_1_3 BL BLB W_1_1_3 W_1_1_3_bar CIM_cell
X4 I11_inv O_1_1_4 WL_1_4 BL BLB W_1_1_4 W_1_1_4_bar CIM_cell
X5 I12_inv O_1_2_1 WL_1_1 BL BLB W_1_2_1 W_1_2_1_bar CIM_cell
X6 I12_inv O_1_2_2 WL_1_2 BL BLB W_1_2_2 W_1_2_2_bar CIM_cell
X7 I12_inv O_1_2_3 WL_1_3 BL BLB W_1_2_3 W_1_2_3_bar CIM_cell
X8 I12_inv O_1_2_4 WL_1_4 BL BLB W_1_2_4 W_1_2_4_bar CIM_cell
X9 I13_inv O_1_3_1 WL_1_1 BL BLB W_1_3_1 W_1_3_1_bar CIM_cell
X10 I13_inv O_1_3_2 WL_1_2 BL BLB W_1_3_2 W_1_3_2_bar CIM_cell
X11 I13_inv O_1_3_3 WL_1_3 BL BLB W_1_3_3 W_1_3_3_bar CIM_cell
X12 I13_inv O_1_3_4 WL_1_4 BL BLB W_1_3_4 W_1_3_4_bar CIM_cell
X13 I14_inv O_1_4_1 WL_1_1 BL BLB W_1_4_1 W_1_4_1_bar CIM_cell
X14 I14_inv O_1_4_2 WL_1_2 BL BLB W_1_4_2 W_1_4_2_bar CIM_cell
X15 I14_inv O_1_4_3 WL_1_3 BL BLB W_1_4_3 W_1_4_3_bar CIM_cell
X16 I14_inv O_1_4_4 WL_1_4 BL BLB W_1_4_4 W_1_4_4_bar CIM_cell
X17 I15_inv O_1_5_1 WL_1_1 BL BLB W_1_5_1 W_1_5_1_bar CIM_cell
X18 I15_inv O_1_5_2 WL_1_2 BL BLB W_1_5_2 W_1_5_2_bar CIM_cell
X19 I15_inv O_1_5_3 WL_1_3 BL BLB W_1_5_3 W_1_5_3_bar CIM_cell
X20 I15_inv O_1_5_4 WL_1_4 BL BLB W_1_5_4 W_1_5_4_bar CIM_cell
X21 I16_inv O_1_6_1 WL_1_1 BL BLB W_1_6_1 W_1_6_1_bar CIM_cell
X22 I16_inv O_1_6_2 WL_1_2 BL BLB W_1_6_2 W_1_6_2_bar CIM_cell
X23 I16_inv O_1_6_3 WL_1_3 BL BLB W_1_6_3 W_1_6_3_bar CIM_cell
X24 I16_inv O_1_6_4 WL_1_4 BL BLB W_1_6_4 W_1_6_4_bar CIM_cell
X25 I17_inv O_1_7_1 WL_1_1 BL BLB W_1_7_1 W_1_7_1_bar CIM_cell
X26 I17_inv O_1_7_2 WL_1_2 BL BLB W_1_7_2 W_1_7_2_bar CIM_cell
X27 I17_inv O_1_7_3 WL_1_3 BL BLB W_1_7_3 W_1_7_3_bar CIM_cell
X28 I17_inv O_1_7_4 WL_1_4 BL BLB W_1_7_4 W_1_7_4_bar CIM_cell
X29 I18_inv O_1_8_1 WL_1_1 BL BLB W_1_8_1 W_1_8_1_bar CIM_cell
X30 I18_inv O_1_8_2 WL_1_2 BL BLB W_1_8_2 W_1_8_2_bar CIM_cell
X31 I18_inv O_1_8_3 WL_1_3 BL BLB W_1_8_3 W_1_8_3_bar CIM_cell
X32 I18_inv O_1_8_4 WL_1_4 BL BLB W_1_8_4 W_1_8_4_bar CIM_cell
X33 I19_inv O_1_9_1 WL_1_1 BL BLB W_1_9_1 W_1_9_1_bar CIM_cell
X34 I19_inv O_1_9_2 WL_1_2 BL BLB W_1_9_2 W_1_9_2_bar CIM_cell
X35 I19_inv O_1_9_3 WL_1_3 BL BLB W_1_9_3 W_1_9_3_bar CIM_cell
X36 I19_inv O_1_9_4 WL_1_4 BL BLB W_1_9_4 W_1_9_4_bar CIM_cell
X37 I110_inv O_1_10_1 WL_1_1 BL BLB W_1_10_1 W_1_10_1_bar CIM_cell
X38 I110_inv O_1_10_2 WL_1_2 BL BLB W_1_10_2 W_1_10_2_bar CIM_cell
X39 I110_inv O_1_10_3 WL_1_3 BL BLB W_1_10_3 W_1_10_3_bar CIM_cell
X40 I110_inv O_1_10_4 WL_1_4 BL BLB W_1_10_4 W_1_10_4_bar CIM_cell
X41 I111_inv O_1_11_1 WL_1_1 BL BLB W_1_11_1 W_1_11_1_bar CIM_cell
X42 I111_inv O_1_11_2 WL_1_2 BL BLB W_1_11_2 W_1_11_2_bar CIM_cell
X43 I111_inv O_1_11_3 WL_1_3 BL BLB W_1_11_3 W_1_11_3_bar CIM_cell
X44 I111_inv O_1_11_4 WL_1_4 BL BLB W_1_11_4 W_1_11_4_bar CIM_cell
X45 I112_inv O_1_12_1 WL_1_1 BL BLB W_1_12_1 W_1_12_1_bar CIM_cell
X46 I112_inv O_1_12_2 WL_1_2 BL BLB W_1_12_2 W_1_12_2_bar CIM_cell
X47 I112_inv O_1_12_3 WL_1_3 BL BLB W_1_12_3 W_1_12_3_bar CIM_cell
X48 I112_inv O_1_12_4 WL_1_4 BL BLB W_1_12_4 W_1_12_4_bar CIM_cell
X49 I113_inv O_1_13_1 WL_1_1 BL BLB W_1_13_1 W_1_13_1_bar CIM_cell
X50 I113_inv O_1_13_2 WL_1_2 BL BLB W_1_13_2 W_1_13_2_bar CIM_cell
X51 I113_inv O_1_13_3 WL_1_3 BL BLB W_1_13_3 W_1_13_3_bar CIM_cell
X52 I113_inv O_1_13_4 WL_1_4 BL BLB W_1_13_4 W_1_13_4_bar CIM_cell
X53 I114_inv O_1_14_1 WL_1_1 BL BLB W_1_14_1 W_1_14_1_bar CIM_cell
X54 I114_inv O_1_14_2 WL_1_2 BL BLB W_1_14_2 W_1_14_2_bar CIM_cell
X55 I114_inv O_1_14_3 WL_1_3 BL BLB W_1_14_3 W_1_14_3_bar CIM_cell
X56 I114_inv O_1_14_4 WL_1_4 BL BLB W_1_14_4 W_1_14_4_bar CIM_cell
X57 I115_inv O_1_15_1 WL_1_1 BL BLB W_1_15_1 W_1_15_1_bar CIM_cell
X58 I115_inv O_1_15_2 WL_1_2 BL BLB W_1_15_2 W_1_15_2_bar CIM_cell
X59 I115_inv O_1_15_3 WL_1_3 BL BLB W_1_15_3 W_1_15_3_bar CIM_cell
X60 I115_inv O_1_15_4 WL_1_4 BL BLB W_1_15_4 W_1_15_4_bar CIM_cell
X61 I116_inv O_1_16_1 WL_1_1 BL BLB W_1_16_1 W_1_16_1_bar CIM_cell
X62 I116_inv O_1_16_2 WL_1_2 BL BLB W_1_16_2 W_1_16_2_bar CIM_cell
X63 I116_inv O_1_16_3 WL_1_3 BL BLB W_1_16_3 W_1_16_3_bar CIM_cell
X64 I116_inv O_1_16_4 WL_1_4 BL BLB W_1_16_4 W_1_16_4_bar CIM_cell
X65 I117_inv O_1_17_1 WL_1_1 BL BLB W_1_17_1 W_1_17_1_bar CIM_cell
X66 I117_inv O_1_17_2 WL_1_2 BL BLB W_1_17_2 W_1_17_2_bar CIM_cell
X67 I117_inv O_1_17_3 WL_1_3 BL BLB W_1_17_3 W_1_17_3_bar CIM_cell
X68 I117_inv O_1_17_4 WL_1_4 BL BLB W_1_17_4 W_1_17_4_bar CIM_cell
X69 I118_inv O_1_18_1 WL_1_1 BL BLB W_1_18_1 W_1_18_1_bar CIM_cell
X70 I118_inv O_1_18_2 WL_1_2 BL BLB W_1_18_2 W_1_18_2_bar CIM_cell
X71 I118_inv O_1_18_3 WL_1_3 BL BLB W_1_18_3 W_1_18_3_bar CIM_cell
X72 I118_inv O_1_18_4 WL_1_4 BL BLB W_1_18_4 W_1_18_4_bar CIM_cell
X73 I119_inv O_1_19_1 WL_1_1 BL BLB W_1_19_1 W_1_19_1_bar CIM_cell
X74 I119_inv O_1_19_2 WL_1_2 BL BLB W_1_19_2 W_1_19_2_bar CIM_cell
X75 I119_inv O_1_19_3 WL_1_3 BL BLB W_1_19_3 W_1_19_3_bar CIM_cell
X76 I119_inv O_1_19_4 WL_1_4 BL BLB W_1_19_4 W_1_19_4_bar CIM_cell
X77 I120_inv O_1_20_1 WL_1_1 BL BLB W_1_20_1 W_1_20_1_bar CIM_cell
X78 I120_inv O_1_20_2 WL_1_2 BL BLB W_1_20_2 W_1_20_2_bar CIM_cell
X79 I120_inv O_1_20_3 WL_1_3 BL BLB W_1_20_3 W_1_20_3_bar CIM_cell
X80 I120_inv O_1_20_4 WL_1_4 BL BLB W_1_20_4 W_1_20_4_bar CIM_cell
X81 I121_inv O_1_21_1 WL_1_1 BL BLB W_1_21_1 W_1_21_1_bar CIM_cell
X82 I121_inv O_1_21_2 WL_1_2 BL BLB W_1_21_2 W_1_21_2_bar CIM_cell
X83 I121_inv O_1_21_3 WL_1_3 BL BLB W_1_21_3 W_1_21_3_bar CIM_cell
X84 I121_inv O_1_21_4 WL_1_4 BL BLB W_1_21_4 W_1_21_4_bar CIM_cell
X85 I122_inv O_1_22_1 WL_1_1 BL BLB W_1_22_1 W_1_22_1_bar CIM_cell
X86 I122_inv O_1_22_2 WL_1_2 BL BLB W_1_22_2 W_1_22_2_bar CIM_cell
X87 I122_inv O_1_22_3 WL_1_3 BL BLB W_1_22_3 W_1_22_3_bar CIM_cell
X88 I122_inv O_1_22_4 WL_1_4 BL BLB W_1_22_4 W_1_22_4_bar CIM_cell
X89 I123_inv O_1_23_1 WL_1_1 BL BLB W_1_23_1 W_1_23_1_bar CIM_cell
X90 I123_inv O_1_23_2 WL_1_2 BL BLB W_1_23_2 W_1_23_2_bar CIM_cell
X91 I123_inv O_1_23_3 WL_1_3 BL BLB W_1_23_3 W_1_23_3_bar CIM_cell
X92 I123_inv O_1_23_4 WL_1_4 BL BLB W_1_23_4 W_1_23_4_bar CIM_cell
X93 I124_inv O_1_24_1 WL_1_1 BL BLB W_1_24_1 W_1_24_1_bar CIM_cell
X94 I124_inv O_1_24_2 WL_1_2 BL BLB W_1_24_2 W_1_24_2_bar CIM_cell
X95 I124_inv O_1_24_3 WL_1_3 BL BLB W_1_24_3 W_1_24_3_bar CIM_cell
X96 I124_inv O_1_24_4 WL_1_4 BL BLB W_1_24_4 W_1_24_4_bar CIM_cell
X97 I125_inv O_1_25_1 WL_1_1 BL BLB W_1_25_1 W_1_25_1_bar CIM_cell
X98 I125_inv O_1_25_2 WL_1_2 BL BLB W_1_25_2 W_1_25_2_bar CIM_cell
X99 I125_inv O_1_25_3 WL_1_3 BL BLB W_1_25_3 W_1_25_3_bar CIM_cell
X100 I125_inv O_1_25_4 WL_1_4 BL BLB W_1_25_4 W_1_25_4_bar CIM_cell
X101 I126_inv O_1_26_1 WL_1_1 BL BLB W_1_26_1 W_1_26_1_bar CIM_cell
X102 I126_inv O_1_26_2 WL_1_2 BL BLB W_1_26_2 W_1_26_2_bar CIM_cell
X103 I126_inv O_1_26_3 WL_1_3 BL BLB W_1_26_3 W_1_26_3_bar CIM_cell
X104 I126_inv O_1_26_4 WL_1_4 BL BLB W_1_26_4 W_1_26_4_bar CIM_cell
X105 I127_inv O_1_27_1 WL_1_1 BL BLB W_1_27_1 W_1_27_1_bar CIM_cell
X106 I127_inv O_1_27_2 WL_1_2 BL BLB W_1_27_2 W_1_27_2_bar CIM_cell
X107 I127_inv O_1_27_3 WL_1_3 BL BLB W_1_27_3 W_1_27_3_bar CIM_cell
X108 I127_inv O_1_27_4 WL_1_4 BL BLB W_1_27_4 W_1_27_4_bar CIM_cell
X109 I128_inv O_1_28_1 WL_1_1 BL BLB W_1_28_1 W_1_28_1_bar CIM_cell
X110 I128_inv O_1_28_2 WL_1_2 BL BLB W_1_28_2 W_1_28_2_bar CIM_cell
X111 I128_inv O_1_28_3 WL_1_3 BL BLB W_1_28_3 W_1_28_3_bar CIM_cell
X112 I128_inv O_1_28_4 WL_1_4 BL BLB W_1_28_4 W_1_28_4_bar CIM_cell
X113 I129_inv O_1_29_1 WL_1_1 BL BLB W_1_29_1 W_1_29_1_bar CIM_cell
X114 I129_inv O_1_29_2 WL_1_2 BL BLB W_1_29_2 W_1_29_2_bar CIM_cell
X115 I129_inv O_1_29_3 WL_1_3 BL BLB W_1_29_3 W_1_29_3_bar CIM_cell
X116 I129_inv O_1_29_4 WL_1_4 BL BLB W_1_29_4 W_1_29_4_bar CIM_cell
X117 I130_inv O_1_30_1 WL_1_1 BL BLB W_1_30_1 W_1_30_1_bar CIM_cell
X118 I130_inv O_1_30_2 WL_1_2 BL BLB W_1_30_2 W_1_30_2_bar CIM_cell
X119 I130_inv O_1_30_3 WL_1_3 BL BLB W_1_30_3 W_1_30_3_bar CIM_cell
X120 I130_inv O_1_30_4 WL_1_4 BL BLB W_1_30_4 W_1_30_4_bar CIM_cell
X121 I131_inv O_1_31_1 WL_1_1 BL BLB W_1_31_1 W_1_31_1_bar CIM_cell
X122 I131_inv O_1_31_2 WL_1_2 BL BLB W_1_31_2 W_1_31_2_bar CIM_cell
X123 I131_inv O_1_31_3 WL_1_3 BL BLB W_1_31_3 W_1_31_3_bar CIM_cell
X124 I131_inv O_1_31_4 WL_1_4 BL BLB W_1_31_4 W_1_31_4_bar CIM_cell
X125 I132_inv O_1_32_1 WL_1_1 BL BLB W_1_32_1 W_1_32_1_bar CIM_cell
X126 I132_inv O_1_32_2 WL_1_2 BL BLB W_1_32_2 W_1_32_2_bar CIM_cell
X127 I132_inv O_1_32_3 WL_1_3 BL BLB W_1_32_3 W_1_32_3_bar CIM_cell
X128 I132_inv O_1_32_4 WL_1_4 BL BLB W_1_32_4 W_1_32_4_bar CIM_cell
X129 I21_inv O_2_1_1 WL_2_1 BL BLB W_2_1_1 W_2_1_1_bar CIM_cell
X130 I21_inv O_2_1_2 WL_2_2 BL BLB W_2_1_2 W_2_1_2_bar CIM_cell
X131 I21_inv O_2_1_3 WL_2_3 BL BLB W_2_1_3 W_2_1_3_bar CIM_cell
X132 I21_inv O_2_1_4 WL_2_4 BL BLB W_2_1_4 W_2_1_4_bar CIM_cell
X133 I22_inv O_2_2_1 WL_2_1 BL BLB W_2_2_1 W_2_2_1_bar CIM_cell
X134 I22_inv O_2_2_2 WL_2_2 BL BLB W_2_2_2 W_2_2_2_bar CIM_cell
X135 I22_inv O_2_2_3 WL_2_3 BL BLB W_2_2_3 W_2_2_3_bar CIM_cell
X136 I22_inv O_2_2_4 WL_2_4 BL BLB W_2_2_4 W_2_2_4_bar CIM_cell
X137 I23_inv O_2_3_1 WL_2_1 BL BLB W_2_3_1 W_2_3_1_bar CIM_cell
X138 I23_inv O_2_3_2 WL_2_2 BL BLB W_2_3_2 W_2_3_2_bar CIM_cell
X139 I23_inv O_2_3_3 WL_2_3 BL BLB W_2_3_3 W_2_3_3_bar CIM_cell
X140 I23_inv O_2_3_4 WL_2_4 BL BLB W_2_3_4 W_2_3_4_bar CIM_cell
X141 I24_inv O_2_4_1 WL_2_1 BL BLB W_2_4_1 W_2_4_1_bar CIM_cell
X142 I24_inv O_2_4_2 WL_2_2 BL BLB W_2_4_2 W_2_4_2_bar CIM_cell
X143 I24_inv O_2_4_3 WL_2_3 BL BLB W_2_4_3 W_2_4_3_bar CIM_cell
X144 I24_inv O_2_4_4 WL_2_4 BL BLB W_2_4_4 W_2_4_4_bar CIM_cell
X145 I25_inv O_2_5_1 WL_2_1 BL BLB W_2_5_1 W_2_5_1_bar CIM_cell
X146 I25_inv O_2_5_2 WL_2_2 BL BLB W_2_5_2 W_2_5_2_bar CIM_cell
X147 I25_inv O_2_5_3 WL_2_3 BL BLB W_2_5_3 W_2_5_3_bar CIM_cell
X148 I25_inv O_2_5_4 WL_2_4 BL BLB W_2_5_4 W_2_5_4_bar CIM_cell
X149 I26_inv O_2_6_1 WL_2_1 BL BLB W_2_6_1 W_2_6_1_bar CIM_cell
X150 I26_inv O_2_6_2 WL_2_2 BL BLB W_2_6_2 W_2_6_2_bar CIM_cell
X151 I26_inv O_2_6_3 WL_2_3 BL BLB W_2_6_3 W_2_6_3_bar CIM_cell
X152 I26_inv O_2_6_4 WL_2_4 BL BLB W_2_6_4 W_2_6_4_bar CIM_cell
X153 I27_inv O_2_7_1 WL_2_1 BL BLB W_2_7_1 W_2_7_1_bar CIM_cell
X154 I27_inv O_2_7_2 WL_2_2 BL BLB W_2_7_2 W_2_7_2_bar CIM_cell
X155 I27_inv O_2_7_3 WL_2_3 BL BLB W_2_7_3 W_2_7_3_bar CIM_cell
X156 I27_inv O_2_7_4 WL_2_4 BL BLB W_2_7_4 W_2_7_4_bar CIM_cell
X157 I28_inv O_2_8_1 WL_2_1 BL BLB W_2_8_1 W_2_8_1_bar CIM_cell
X158 I28_inv O_2_8_2 WL_2_2 BL BLB W_2_8_2 W_2_8_2_bar CIM_cell
X159 I28_inv O_2_8_3 WL_2_3 BL BLB W_2_8_3 W_2_8_3_bar CIM_cell
X160 I28_inv O_2_8_4 WL_2_4 BL BLB W_2_8_4 W_2_8_4_bar CIM_cell
X161 I29_inv O_2_9_1 WL_2_1 BL BLB W_2_9_1 W_2_9_1_bar CIM_cell
X162 I29_inv O_2_9_2 WL_2_2 BL BLB W_2_9_2 W_2_9_2_bar CIM_cell
X163 I29_inv O_2_9_3 WL_2_3 BL BLB W_2_9_3 W_2_9_3_bar CIM_cell
X164 I29_inv O_2_9_4 WL_2_4 BL BLB W_2_9_4 W_2_9_4_bar CIM_cell
X165 I210_inv O_2_10_1 WL_2_1 BL BLB W_2_10_1 W_2_10_1_bar CIM_cell
X166 I210_inv O_2_10_2 WL_2_2 BL BLB W_2_10_2 W_2_10_2_bar CIM_cell
X167 I210_inv O_2_10_3 WL_2_3 BL BLB W_2_10_3 W_2_10_3_bar CIM_cell
X168 I210_inv O_2_10_4 WL_2_4 BL BLB W_2_10_4 W_2_10_4_bar CIM_cell
X169 I211_inv O_2_11_1 WL_2_1 BL BLB W_2_11_1 W_2_11_1_bar CIM_cell
X170 I211_inv O_2_11_2 WL_2_2 BL BLB W_2_11_2 W_2_11_2_bar CIM_cell
X171 I211_inv O_2_11_3 WL_2_3 BL BLB W_2_11_3 W_2_11_3_bar CIM_cell
X172 I211_inv O_2_11_4 WL_2_4 BL BLB W_2_11_4 W_2_11_4_bar CIM_cell
X173 I212_inv O_2_12_1 WL_2_1 BL BLB W_2_12_1 W_2_12_1_bar CIM_cell
X174 I212_inv O_2_12_2 WL_2_2 BL BLB W_2_12_2 W_2_12_2_bar CIM_cell
X175 I212_inv O_2_12_3 WL_2_3 BL BLB W_2_12_3 W_2_12_3_bar CIM_cell
X176 I212_inv O_2_12_4 WL_2_4 BL BLB W_2_12_4 W_2_12_4_bar CIM_cell
X177 I213_inv O_2_13_1 WL_2_1 BL BLB W_2_13_1 W_2_13_1_bar CIM_cell
X178 I213_inv O_2_13_2 WL_2_2 BL BLB W_2_13_2 W_2_13_2_bar CIM_cell
X179 I213_inv O_2_13_3 WL_2_3 BL BLB W_2_13_3 W_2_13_3_bar CIM_cell
X180 I213_inv O_2_13_4 WL_2_4 BL BLB W_2_13_4 W_2_13_4_bar CIM_cell
X181 I214_inv O_2_14_1 WL_2_1 BL BLB W_2_14_1 W_2_14_1_bar CIM_cell
X182 I214_inv O_2_14_2 WL_2_2 BL BLB W_2_14_2 W_2_14_2_bar CIM_cell
X183 I214_inv O_2_14_3 WL_2_3 BL BLB W_2_14_3 W_2_14_3_bar CIM_cell
X184 I214_inv O_2_14_4 WL_2_4 BL BLB W_2_14_4 W_2_14_4_bar CIM_cell
X185 I215_inv O_2_15_1 WL_2_1 BL BLB W_2_15_1 W_2_15_1_bar CIM_cell
X186 I215_inv O_2_15_2 WL_2_2 BL BLB W_2_15_2 W_2_15_2_bar CIM_cell
X187 I215_inv O_2_15_3 WL_2_3 BL BLB W_2_15_3 W_2_15_3_bar CIM_cell
X188 I215_inv O_2_15_4 WL_2_4 BL BLB W_2_15_4 W_2_15_4_bar CIM_cell
X189 I216_inv O_2_16_1 WL_2_1 BL BLB W_2_16_1 W_2_16_1_bar CIM_cell
X190 I216_inv O_2_16_2 WL_2_2 BL BLB W_2_16_2 W_2_16_2_bar CIM_cell
X191 I216_inv O_2_16_3 WL_2_3 BL BLB W_2_16_3 W_2_16_3_bar CIM_cell
X192 I216_inv O_2_16_4 WL_2_4 BL BLB W_2_16_4 W_2_16_4_bar CIM_cell
X193 I217_inv O_2_17_1 WL_2_1 BL BLB W_2_17_1 W_2_17_1_bar CIM_cell
X194 I217_inv O_2_17_2 WL_2_2 BL BLB W_2_17_2 W_2_17_2_bar CIM_cell
X195 I217_inv O_2_17_3 WL_2_3 BL BLB W_2_17_3 W_2_17_3_bar CIM_cell
X196 I217_inv O_2_17_4 WL_2_4 BL BLB W_2_17_4 W_2_17_4_bar CIM_cell
X197 I218_inv O_2_18_1 WL_2_1 BL BLB W_2_18_1 W_2_18_1_bar CIM_cell
X198 I218_inv O_2_18_2 WL_2_2 BL BLB W_2_18_2 W_2_18_2_bar CIM_cell
X199 I218_inv O_2_18_3 WL_2_3 BL BLB W_2_18_3 W_2_18_3_bar CIM_cell
X200 I218_inv O_2_18_4 WL_2_4 BL BLB W_2_18_4 W_2_18_4_bar CIM_cell
X201 I219_inv O_2_19_1 WL_2_1 BL BLB W_2_19_1 W_2_19_1_bar CIM_cell
X202 I219_inv O_2_19_2 WL_2_2 BL BLB W_2_19_2 W_2_19_2_bar CIM_cell
X203 I219_inv O_2_19_3 WL_2_3 BL BLB W_2_19_3 W_2_19_3_bar CIM_cell
X204 I219_inv O_2_19_4 WL_2_4 BL BLB W_2_19_4 W_2_19_4_bar CIM_cell
X205 I220_inv O_2_20_1 WL_2_1 BL BLB W_2_20_1 W_2_20_1_bar CIM_cell
X206 I220_inv O_2_20_2 WL_2_2 BL BLB W_2_20_2 W_2_20_2_bar CIM_cell
X207 I220_inv O_2_20_3 WL_2_3 BL BLB W_2_20_3 W_2_20_3_bar CIM_cell
X208 I220_inv O_2_20_4 WL_2_4 BL BLB W_2_20_4 W_2_20_4_bar CIM_cell
X209 I221_inv O_2_21_1 WL_2_1 BL BLB W_2_21_1 W_2_21_1_bar CIM_cell
X210 I221_inv O_2_21_2 WL_2_2 BL BLB W_2_21_2 W_2_21_2_bar CIM_cell
X211 I221_inv O_2_21_3 WL_2_3 BL BLB W_2_21_3 W_2_21_3_bar CIM_cell
X212 I221_inv O_2_21_4 WL_2_4 BL BLB W_2_21_4 W_2_21_4_bar CIM_cell
X213 I222_inv O_2_22_1 WL_2_1 BL BLB W_2_22_1 W_2_22_1_bar CIM_cell
X214 I222_inv O_2_22_2 WL_2_2 BL BLB W_2_22_2 W_2_22_2_bar CIM_cell
X215 I222_inv O_2_22_3 WL_2_3 BL BLB W_2_22_3 W_2_22_3_bar CIM_cell
X216 I222_inv O_2_22_4 WL_2_4 BL BLB W_2_22_4 W_2_22_4_bar CIM_cell
X217 I223_inv O_2_23_1 WL_2_1 BL BLB W_2_23_1 W_2_23_1_bar CIM_cell
X218 I223_inv O_2_23_2 WL_2_2 BL BLB W_2_23_2 W_2_23_2_bar CIM_cell
X219 I223_inv O_2_23_3 WL_2_3 BL BLB W_2_23_3 W_2_23_3_bar CIM_cell
X220 I223_inv O_2_23_4 WL_2_4 BL BLB W_2_23_4 W_2_23_4_bar CIM_cell
X221 I224_inv O_2_24_1 WL_2_1 BL BLB W_2_24_1 W_2_24_1_bar CIM_cell
X222 I224_inv O_2_24_2 WL_2_2 BL BLB W_2_24_2 W_2_24_2_bar CIM_cell
X223 I224_inv O_2_24_3 WL_2_3 BL BLB W_2_24_3 W_2_24_3_bar CIM_cell
X224 I224_inv O_2_24_4 WL_2_4 BL BLB W_2_24_4 W_2_24_4_bar CIM_cell
X225 I225_inv O_2_25_1 WL_2_1 BL BLB W_2_25_1 W_2_25_1_bar CIM_cell
X226 I225_inv O_2_25_2 WL_2_2 BL BLB W_2_25_2 W_2_25_2_bar CIM_cell
X227 I225_inv O_2_25_3 WL_2_3 BL BLB W_2_25_3 W_2_25_3_bar CIM_cell
X228 I225_inv O_2_25_4 WL_2_4 BL BLB W_2_25_4 W_2_25_4_bar CIM_cell
X229 I226_inv O_2_26_1 WL_2_1 BL BLB W_2_26_1 W_2_26_1_bar CIM_cell
X230 I226_inv O_2_26_2 WL_2_2 BL BLB W_2_26_2 W_2_26_2_bar CIM_cell
X231 I226_inv O_2_26_3 WL_2_3 BL BLB W_2_26_3 W_2_26_3_bar CIM_cell
X232 I226_inv O_2_26_4 WL_2_4 BL BLB W_2_26_4 W_2_26_4_bar CIM_cell
X233 I227_inv O_2_27_1 WL_2_1 BL BLB W_2_27_1 W_2_27_1_bar CIM_cell
X234 I227_inv O_2_27_2 WL_2_2 BL BLB W_2_27_2 W_2_27_2_bar CIM_cell
X235 I227_inv O_2_27_3 WL_2_3 BL BLB W_2_27_3 W_2_27_3_bar CIM_cell
X236 I227_inv O_2_27_4 WL_2_4 BL BLB W_2_27_4 W_2_27_4_bar CIM_cell
X237 I228_inv O_2_28_1 WL_2_1 BL BLB W_2_28_1 W_2_28_1_bar CIM_cell
X238 I228_inv O_2_28_2 WL_2_2 BL BLB W_2_28_2 W_2_28_2_bar CIM_cell
X239 I228_inv O_2_28_3 WL_2_3 BL BLB W_2_28_3 W_2_28_3_bar CIM_cell
X240 I228_inv O_2_28_4 WL_2_4 BL BLB W_2_28_4 W_2_28_4_bar CIM_cell
X241 I229_inv O_2_29_1 WL_2_1 BL BLB W_2_29_1 W_2_29_1_bar CIM_cell
X242 I229_inv O_2_29_2 WL_2_2 BL BLB W_2_29_2 W_2_29_2_bar CIM_cell
X243 I229_inv O_2_29_3 WL_2_3 BL BLB W_2_29_3 W_2_29_3_bar CIM_cell
X244 I229_inv O_2_29_4 WL_2_4 BL BLB W_2_29_4 W_2_29_4_bar CIM_cell
X245 I230_inv O_2_30_1 WL_2_1 BL BLB W_2_30_1 W_2_30_1_bar CIM_cell
X246 I230_inv O_2_30_2 WL_2_2 BL BLB W_2_30_2 W_2_30_2_bar CIM_cell
X247 I230_inv O_2_30_3 WL_2_3 BL BLB W_2_30_3 W_2_30_3_bar CIM_cell
X248 I230_inv O_2_30_4 WL_2_4 BL BLB W_2_30_4 W_2_30_4_bar CIM_cell
X249 I231_inv O_2_31_1 WL_2_1 BL BLB W_2_31_1 W_2_31_1_bar CIM_cell
X250 I231_inv O_2_31_2 WL_2_2 BL BLB W_2_31_2 W_2_31_2_bar CIM_cell
X251 I231_inv O_2_31_3 WL_2_3 BL BLB W_2_31_3 W_2_31_3_bar CIM_cell
X252 I231_inv O_2_31_4 WL_2_4 BL BLB W_2_31_4 W_2_31_4_bar CIM_cell
X253 I232_inv O_2_32_1 WL_2_1 BL BLB W_2_32_1 W_2_32_1_bar CIM_cell
X254 I232_inv O_2_32_2 WL_2_2 BL BLB W_2_32_2 W_2_32_2_bar CIM_cell
X255 I232_inv O_2_32_3 WL_2_3 BL BLB W_2_32_3 W_2_32_3_bar CIM_cell
X256 I232_inv O_2_32_4 WL_2_4 BL BLB W_2_32_4 W_2_32_4_bar CIM_cell
X257 I31_inv O_3_1_1 WL_3_1 BL BLB W_3_1_1 W_3_1_1_bar CIM_cell
X258 I31_inv O_3_1_2 WL_3_2 BL BLB W_3_1_2 W_3_1_2_bar CIM_cell
X259 I31_inv O_3_1_3 WL_3_3 BL BLB W_3_1_3 W_3_1_3_bar CIM_cell
X260 I31_inv O_3_1_4 WL_3_4 BL BLB W_3_1_4 W_3_1_4_bar CIM_cell
X261 I32_inv O_3_2_1 WL_3_1 BL BLB W_3_2_1 W_3_2_1_bar CIM_cell
X262 I32_inv O_3_2_2 WL_3_2 BL BLB W_3_2_2 W_3_2_2_bar CIM_cell
X263 I32_inv O_3_2_3 WL_3_3 BL BLB W_3_2_3 W_3_2_3_bar CIM_cell
X264 I32_inv O_3_2_4 WL_3_4 BL BLB W_3_2_4 W_3_2_4_bar CIM_cell
X265 I33_inv O_3_3_1 WL_3_1 BL BLB W_3_3_1 W_3_3_1_bar CIM_cell
X266 I33_inv O_3_3_2 WL_3_2 BL BLB W_3_3_2 W_3_3_2_bar CIM_cell
X267 I33_inv O_3_3_3 WL_3_3 BL BLB W_3_3_3 W_3_3_3_bar CIM_cell
X268 I33_inv O_3_3_4 WL_3_4 BL BLB W_3_3_4 W_3_3_4_bar CIM_cell
X269 I34_inv O_3_4_1 WL_3_1 BL BLB W_3_4_1 W_3_4_1_bar CIM_cell
X270 I34_inv O_3_4_2 WL_3_2 BL BLB W_3_4_2 W_3_4_2_bar CIM_cell
X271 I34_inv O_3_4_3 WL_3_3 BL BLB W_3_4_3 W_3_4_3_bar CIM_cell
X272 I34_inv O_3_4_4 WL_3_4 BL BLB W_3_4_4 W_3_4_4_bar CIM_cell
X273 I35_inv O_3_5_1 WL_3_1 BL BLB W_3_5_1 W_3_5_1_bar CIM_cell
X274 I35_inv O_3_5_2 WL_3_2 BL BLB W_3_5_2 W_3_5_2_bar CIM_cell
X275 I35_inv O_3_5_3 WL_3_3 BL BLB W_3_5_3 W_3_5_3_bar CIM_cell
X276 I35_inv O_3_5_4 WL_3_4 BL BLB W_3_5_4 W_3_5_4_bar CIM_cell
X277 I36_inv O_3_6_1 WL_3_1 BL BLB W_3_6_1 W_3_6_1_bar CIM_cell
X278 I36_inv O_3_6_2 WL_3_2 BL BLB W_3_6_2 W_3_6_2_bar CIM_cell
X279 I36_inv O_3_6_3 WL_3_3 BL BLB W_3_6_3 W_3_6_3_bar CIM_cell
X280 I36_inv O_3_6_4 WL_3_4 BL BLB W_3_6_4 W_3_6_4_bar CIM_cell
X281 I37_inv O_3_7_1 WL_3_1 BL BLB W_3_7_1 W_3_7_1_bar CIM_cell
X282 I37_inv O_3_7_2 WL_3_2 BL BLB W_3_7_2 W_3_7_2_bar CIM_cell
X283 I37_inv O_3_7_3 WL_3_3 BL BLB W_3_7_3 W_3_7_3_bar CIM_cell
X284 I37_inv O_3_7_4 WL_3_4 BL BLB W_3_7_4 W_3_7_4_bar CIM_cell
X285 I38_inv O_3_8_1 WL_3_1 BL BLB W_3_8_1 W_3_8_1_bar CIM_cell
X286 I38_inv O_3_8_2 WL_3_2 BL BLB W_3_8_2 W_3_8_2_bar CIM_cell
X287 I38_inv O_3_8_3 WL_3_3 BL BLB W_3_8_3 W_3_8_3_bar CIM_cell
X288 I38_inv O_3_8_4 WL_3_4 BL BLB W_3_8_4 W_3_8_4_bar CIM_cell
X289 I39_inv O_3_9_1 WL_3_1 BL BLB W_3_9_1 W_3_9_1_bar CIM_cell
X290 I39_inv O_3_9_2 WL_3_2 BL BLB W_3_9_2 W_3_9_2_bar CIM_cell
X291 I39_inv O_3_9_3 WL_3_3 BL BLB W_3_9_3 W_3_9_3_bar CIM_cell
X292 I39_inv O_3_9_4 WL_3_4 BL BLB W_3_9_4 W_3_9_4_bar CIM_cell
X293 I310_inv O_3_10_1 WL_3_1 BL BLB W_3_10_1 W_3_10_1_bar CIM_cell
X294 I310_inv O_3_10_2 WL_3_2 BL BLB W_3_10_2 W_3_10_2_bar CIM_cell
X295 I310_inv O_3_10_3 WL_3_3 BL BLB W_3_10_3 W_3_10_3_bar CIM_cell
X296 I310_inv O_3_10_4 WL_3_4 BL BLB W_3_10_4 W_3_10_4_bar CIM_cell
X297 I311_inv O_3_11_1 WL_3_1 BL BLB W_3_11_1 W_3_11_1_bar CIM_cell
X298 I311_inv O_3_11_2 WL_3_2 BL BLB W_3_11_2 W_3_11_2_bar CIM_cell
X299 I311_inv O_3_11_3 WL_3_3 BL BLB W_3_11_3 W_3_11_3_bar CIM_cell
X300 I311_inv O_3_11_4 WL_3_4 BL BLB W_3_11_4 W_3_11_4_bar CIM_cell
X301 I312_inv O_3_12_1 WL_3_1 BL BLB W_3_12_1 W_3_12_1_bar CIM_cell
X302 I312_inv O_3_12_2 WL_3_2 BL BLB W_3_12_2 W_3_12_2_bar CIM_cell
X303 I312_inv O_3_12_3 WL_3_3 BL BLB W_3_12_3 W_3_12_3_bar CIM_cell
X304 I312_inv O_3_12_4 WL_3_4 BL BLB W_3_12_4 W_3_12_4_bar CIM_cell
X305 I313_inv O_3_13_1 WL_3_1 BL BLB W_3_13_1 W_3_13_1_bar CIM_cell
X306 I313_inv O_3_13_2 WL_3_2 BL BLB W_3_13_2 W_3_13_2_bar CIM_cell
X307 I313_inv O_3_13_3 WL_3_3 BL BLB W_3_13_3 W_3_13_3_bar CIM_cell
X308 I313_inv O_3_13_4 WL_3_4 BL BLB W_3_13_4 W_3_13_4_bar CIM_cell
X309 I314_inv O_3_14_1 WL_3_1 BL BLB W_3_14_1 W_3_14_1_bar CIM_cell
X310 I314_inv O_3_14_2 WL_3_2 BL BLB W_3_14_2 W_3_14_2_bar CIM_cell
X311 I314_inv O_3_14_3 WL_3_3 BL BLB W_3_14_3 W_3_14_3_bar CIM_cell
X312 I314_inv O_3_14_4 WL_3_4 BL BLB W_3_14_4 W_3_14_4_bar CIM_cell
X313 I315_inv O_3_15_1 WL_3_1 BL BLB W_3_15_1 W_3_15_1_bar CIM_cell
X314 I315_inv O_3_15_2 WL_3_2 BL BLB W_3_15_2 W_3_15_2_bar CIM_cell
X315 I315_inv O_3_15_3 WL_3_3 BL BLB W_3_15_3 W_3_15_3_bar CIM_cell
X316 I315_inv O_3_15_4 WL_3_4 BL BLB W_3_15_4 W_3_15_4_bar CIM_cell
X317 I316_inv O_3_16_1 WL_3_1 BL BLB W_3_16_1 W_3_16_1_bar CIM_cell
X318 I316_inv O_3_16_2 WL_3_2 BL BLB W_3_16_2 W_3_16_2_bar CIM_cell
X319 I316_inv O_3_16_3 WL_3_3 BL BLB W_3_16_3 W_3_16_3_bar CIM_cell
X320 I316_inv O_3_16_4 WL_3_4 BL BLB W_3_16_4 W_3_16_4_bar CIM_cell
X321 I317_inv O_3_17_1 WL_3_1 BL BLB W_3_17_1 W_3_17_1_bar CIM_cell
X322 I317_inv O_3_17_2 WL_3_2 BL BLB W_3_17_2 W_3_17_2_bar CIM_cell
X323 I317_inv O_3_17_3 WL_3_3 BL BLB W_3_17_3 W_3_17_3_bar CIM_cell
X324 I317_inv O_3_17_4 WL_3_4 BL BLB W_3_17_4 W_3_17_4_bar CIM_cell
X325 I318_inv O_3_18_1 WL_3_1 BL BLB W_3_18_1 W_3_18_1_bar CIM_cell
X326 I318_inv O_3_18_2 WL_3_2 BL BLB W_3_18_2 W_3_18_2_bar CIM_cell
X327 I318_inv O_3_18_3 WL_3_3 BL BLB W_3_18_3 W_3_18_3_bar CIM_cell
X328 I318_inv O_3_18_4 WL_3_4 BL BLB W_3_18_4 W_3_18_4_bar CIM_cell
X329 I319_inv O_3_19_1 WL_3_1 BL BLB W_3_19_1 W_3_19_1_bar CIM_cell
X330 I319_inv O_3_19_2 WL_3_2 BL BLB W_3_19_2 W_3_19_2_bar CIM_cell
X331 I319_inv O_3_19_3 WL_3_3 BL BLB W_3_19_3 W_3_19_3_bar CIM_cell
X332 I319_inv O_3_19_4 WL_3_4 BL BLB W_3_19_4 W_3_19_4_bar CIM_cell
X333 I320_inv O_3_20_1 WL_3_1 BL BLB W_3_20_1 W_3_20_1_bar CIM_cell
X334 I320_inv O_3_20_2 WL_3_2 BL BLB W_3_20_2 W_3_20_2_bar CIM_cell
X335 I320_inv O_3_20_3 WL_3_3 BL BLB W_3_20_3 W_3_20_3_bar CIM_cell
X336 I320_inv O_3_20_4 WL_3_4 BL BLB W_3_20_4 W_3_20_4_bar CIM_cell
X337 I321_inv O_3_21_1 WL_3_1 BL BLB W_3_21_1 W_3_21_1_bar CIM_cell
X338 I321_inv O_3_21_2 WL_3_2 BL BLB W_3_21_2 W_3_21_2_bar CIM_cell
X339 I321_inv O_3_21_3 WL_3_3 BL BLB W_3_21_3 W_3_21_3_bar CIM_cell
X340 I321_inv O_3_21_4 WL_3_4 BL BLB W_3_21_4 W_3_21_4_bar CIM_cell
X341 I322_inv O_3_22_1 WL_3_1 BL BLB W_3_22_1 W_3_22_1_bar CIM_cell
X342 I322_inv O_3_22_2 WL_3_2 BL BLB W_3_22_2 W_3_22_2_bar CIM_cell
X343 I322_inv O_3_22_3 WL_3_3 BL BLB W_3_22_3 W_3_22_3_bar CIM_cell
X344 I322_inv O_3_22_4 WL_3_4 BL BLB W_3_22_4 W_3_22_4_bar CIM_cell
X345 I323_inv O_3_23_1 WL_3_1 BL BLB W_3_23_1 W_3_23_1_bar CIM_cell
X346 I323_inv O_3_23_2 WL_3_2 BL BLB W_3_23_2 W_3_23_2_bar CIM_cell
X347 I323_inv O_3_23_3 WL_3_3 BL BLB W_3_23_3 W_3_23_3_bar CIM_cell
X348 I323_inv O_3_23_4 WL_3_4 BL BLB W_3_23_4 W_3_23_4_bar CIM_cell
X349 I324_inv O_3_24_1 WL_3_1 BL BLB W_3_24_1 W_3_24_1_bar CIM_cell
X350 I324_inv O_3_24_2 WL_3_2 BL BLB W_3_24_2 W_3_24_2_bar CIM_cell
X351 I324_inv O_3_24_3 WL_3_3 BL BLB W_3_24_3 W_3_24_3_bar CIM_cell
X352 I324_inv O_3_24_4 WL_3_4 BL BLB W_3_24_4 W_3_24_4_bar CIM_cell
X353 I325_inv O_3_25_1 WL_3_1 BL BLB W_3_25_1 W_3_25_1_bar CIM_cell
X354 I325_inv O_3_25_2 WL_3_2 BL BLB W_3_25_2 W_3_25_2_bar CIM_cell
X355 I325_inv O_3_25_3 WL_3_3 BL BLB W_3_25_3 W_3_25_3_bar CIM_cell
X356 I325_inv O_3_25_4 WL_3_4 BL BLB W_3_25_4 W_3_25_4_bar CIM_cell
X357 I326_inv O_3_26_1 WL_3_1 BL BLB W_3_26_1 W_3_26_1_bar CIM_cell
X358 I326_inv O_3_26_2 WL_3_2 BL BLB W_3_26_2 W_3_26_2_bar CIM_cell
X359 I326_inv O_3_26_3 WL_3_3 BL BLB W_3_26_3 W_3_26_3_bar CIM_cell
X360 I326_inv O_3_26_4 WL_3_4 BL BLB W_3_26_4 W_3_26_4_bar CIM_cell
X361 I327_inv O_3_27_1 WL_3_1 BL BLB W_3_27_1 W_3_27_1_bar CIM_cell
X362 I327_inv O_3_27_2 WL_3_2 BL BLB W_3_27_2 W_3_27_2_bar CIM_cell
X363 I327_inv O_3_27_3 WL_3_3 BL BLB W_3_27_3 W_3_27_3_bar CIM_cell
X364 I327_inv O_3_27_4 WL_3_4 BL BLB W_3_27_4 W_3_27_4_bar CIM_cell
X365 I328_inv O_3_28_1 WL_3_1 BL BLB W_3_28_1 W_3_28_1_bar CIM_cell
X366 I328_inv O_3_28_2 WL_3_2 BL BLB W_3_28_2 W_3_28_2_bar CIM_cell
X367 I328_inv O_3_28_3 WL_3_3 BL BLB W_3_28_3 W_3_28_3_bar CIM_cell
X368 I328_inv O_3_28_4 WL_3_4 BL BLB W_3_28_4 W_3_28_4_bar CIM_cell
X369 I329_inv O_3_29_1 WL_3_1 BL BLB W_3_29_1 W_3_29_1_bar CIM_cell
X370 I329_inv O_3_29_2 WL_3_2 BL BLB W_3_29_2 W_3_29_2_bar CIM_cell
X371 I329_inv O_3_29_3 WL_3_3 BL BLB W_3_29_3 W_3_29_3_bar CIM_cell
X372 I329_inv O_3_29_4 WL_3_4 BL BLB W_3_29_4 W_3_29_4_bar CIM_cell
X373 I330_inv O_3_30_1 WL_3_1 BL BLB W_3_30_1 W_3_30_1_bar CIM_cell
X374 I330_inv O_3_30_2 WL_3_2 BL BLB W_3_30_2 W_3_30_2_bar CIM_cell
X375 I330_inv O_3_30_3 WL_3_3 BL BLB W_3_30_3 W_3_30_3_bar CIM_cell
X376 I330_inv O_3_30_4 WL_3_4 BL BLB W_3_30_4 W_3_30_4_bar CIM_cell
X377 I331_inv O_3_31_1 WL_3_1 BL BLB W_3_31_1 W_3_31_1_bar CIM_cell
X378 I331_inv O_3_31_2 WL_3_2 BL BLB W_3_31_2 W_3_31_2_bar CIM_cell
X379 I331_inv O_3_31_3 WL_3_3 BL BLB W_3_31_3 W_3_31_3_bar CIM_cell
X380 I331_inv O_3_31_4 WL_3_4 BL BLB W_3_31_4 W_3_31_4_bar CIM_cell
X381 I332_inv O_3_32_1 WL_3_1 BL BLB W_3_32_1 W_3_32_1_bar CIM_cell
X382 I332_inv O_3_32_2 WL_3_2 BL BLB W_3_32_2 W_3_32_2_bar CIM_cell
X383 I332_inv O_3_32_3 WL_3_3 BL BLB W_3_32_3 W_3_32_3_bar CIM_cell
X384 I332_inv O_3_32_4 WL_3_4 BL BLB W_3_32_4 W_3_32_4_bar CIM_cell
X385 I41_inv O_4_1_1 WL_4_1 BL BLB W_4_1_1 W_4_1_1_bar CIM_cell
X386 I41_inv O_4_1_2 WL_4_2 BL BLB W_4_1_2 W_4_1_2_bar CIM_cell
X387 I41_inv O_4_1_3 WL_4_3 BL BLB W_4_1_3 W_4_1_3_bar CIM_cell
X388 I41_inv O_4_1_4 WL_4_4 BL BLB W_4_1_4 W_4_1_4_bar CIM_cell
X389 I42_inv O_4_2_1 WL_4_1 BL BLB W_4_2_1 W_4_2_1_bar CIM_cell
X390 I42_inv O_4_2_2 WL_4_2 BL BLB W_4_2_2 W_4_2_2_bar CIM_cell
X391 I42_inv O_4_2_3 WL_4_3 BL BLB W_4_2_3 W_4_2_3_bar CIM_cell
X392 I42_inv O_4_2_4 WL_4_4 BL BLB W_4_2_4 W_4_2_4_bar CIM_cell
X393 I43_inv O_4_3_1 WL_4_1 BL BLB W_4_3_1 W_4_3_1_bar CIM_cell
X394 I43_inv O_4_3_2 WL_4_2 BL BLB W_4_3_2 W_4_3_2_bar CIM_cell
X395 I43_inv O_4_3_3 WL_4_3 BL BLB W_4_3_3 W_4_3_3_bar CIM_cell
X396 I43_inv O_4_3_4 WL_4_4 BL BLB W_4_3_4 W_4_3_4_bar CIM_cell
X397 I44_inv O_4_4_1 WL_4_1 BL BLB W_4_4_1 W_4_4_1_bar CIM_cell
X398 I44_inv O_4_4_2 WL_4_2 BL BLB W_4_4_2 W_4_4_2_bar CIM_cell
X399 I44_inv O_4_4_3 WL_4_3 BL BLB W_4_4_3 W_4_4_3_bar CIM_cell
X400 I44_inv O_4_4_4 WL_4_4 BL BLB W_4_4_4 W_4_4_4_bar CIM_cell
X401 I45_inv O_4_5_1 WL_4_1 BL BLB W_4_5_1 W_4_5_1_bar CIM_cell
X402 I45_inv O_4_5_2 WL_4_2 BL BLB W_4_5_2 W_4_5_2_bar CIM_cell
X403 I45_inv O_4_5_3 WL_4_3 BL BLB W_4_5_3 W_4_5_3_bar CIM_cell
X404 I45_inv O_4_5_4 WL_4_4 BL BLB W_4_5_4 W_4_5_4_bar CIM_cell
X405 I46_inv O_4_6_1 WL_4_1 BL BLB W_4_6_1 W_4_6_1_bar CIM_cell
X406 I46_inv O_4_6_2 WL_4_2 BL BLB W_4_6_2 W_4_6_2_bar CIM_cell
X407 I46_inv O_4_6_3 WL_4_3 BL BLB W_4_6_3 W_4_6_3_bar CIM_cell
X408 I46_inv O_4_6_4 WL_4_4 BL BLB W_4_6_4 W_4_6_4_bar CIM_cell
X409 I47_inv O_4_7_1 WL_4_1 BL BLB W_4_7_1 W_4_7_1_bar CIM_cell
X410 I47_inv O_4_7_2 WL_4_2 BL BLB W_4_7_2 W_4_7_2_bar CIM_cell
X411 I47_inv O_4_7_3 WL_4_3 BL BLB W_4_7_3 W_4_7_3_bar CIM_cell
X412 I47_inv O_4_7_4 WL_4_4 BL BLB W_4_7_4 W_4_7_4_bar CIM_cell
X413 I48_inv O_4_8_1 WL_4_1 BL BLB W_4_8_1 W_4_8_1_bar CIM_cell
X414 I48_inv O_4_8_2 WL_4_2 BL BLB W_4_8_2 W_4_8_2_bar CIM_cell
X415 I48_inv O_4_8_3 WL_4_3 BL BLB W_4_8_3 W_4_8_3_bar CIM_cell
X416 I48_inv O_4_8_4 WL_4_4 BL BLB W_4_8_4 W_4_8_4_bar CIM_cell
X417 I49_inv O_4_9_1 WL_4_1 BL BLB W_4_9_1 W_4_9_1_bar CIM_cell
X418 I49_inv O_4_9_2 WL_4_2 BL BLB W_4_9_2 W_4_9_2_bar CIM_cell
X419 I49_inv O_4_9_3 WL_4_3 BL BLB W_4_9_3 W_4_9_3_bar CIM_cell
X420 I49_inv O_4_9_4 WL_4_4 BL BLB W_4_9_4 W_4_9_4_bar CIM_cell
X421 I410_inv O_4_10_1 WL_4_1 BL BLB W_4_10_1 W_4_10_1_bar CIM_cell
X422 I410_inv O_4_10_2 WL_4_2 BL BLB W_4_10_2 W_4_10_2_bar CIM_cell
X423 I410_inv O_4_10_3 WL_4_3 BL BLB W_4_10_3 W_4_10_3_bar CIM_cell
X424 I410_inv O_4_10_4 WL_4_4 BL BLB W_4_10_4 W_4_10_4_bar CIM_cell
X425 I411_inv O_4_11_1 WL_4_1 BL BLB W_4_11_1 W_4_11_1_bar CIM_cell
X426 I411_inv O_4_11_2 WL_4_2 BL BLB W_4_11_2 W_4_11_2_bar CIM_cell
X427 I411_inv O_4_11_3 WL_4_3 BL BLB W_4_11_3 W_4_11_3_bar CIM_cell
X428 I411_inv O_4_11_4 WL_4_4 BL BLB W_4_11_4 W_4_11_4_bar CIM_cell
X429 I412_inv O_4_12_1 WL_4_1 BL BLB W_4_12_1 W_4_12_1_bar CIM_cell
X430 I412_inv O_4_12_2 WL_4_2 BL BLB W_4_12_2 W_4_12_2_bar CIM_cell
X431 I412_inv O_4_12_3 WL_4_3 BL BLB W_4_12_3 W_4_12_3_bar CIM_cell
X432 I412_inv O_4_12_4 WL_4_4 BL BLB W_4_12_4 W_4_12_4_bar CIM_cell
X433 I413_inv O_4_13_1 WL_4_1 BL BLB W_4_13_1 W_4_13_1_bar CIM_cell
X434 I413_inv O_4_13_2 WL_4_2 BL BLB W_4_13_2 W_4_13_2_bar CIM_cell
X435 I413_inv O_4_13_3 WL_4_3 BL BLB W_4_13_3 W_4_13_3_bar CIM_cell
X436 I413_inv O_4_13_4 WL_4_4 BL BLB W_4_13_4 W_4_13_4_bar CIM_cell
X437 I414_inv O_4_14_1 WL_4_1 BL BLB W_4_14_1 W_4_14_1_bar CIM_cell
X438 I414_inv O_4_14_2 WL_4_2 BL BLB W_4_14_2 W_4_14_2_bar CIM_cell
X439 I414_inv O_4_14_3 WL_4_3 BL BLB W_4_14_3 W_4_14_3_bar CIM_cell
X440 I414_inv O_4_14_4 WL_4_4 BL BLB W_4_14_4 W_4_14_4_bar CIM_cell
X441 I415_inv O_4_15_1 WL_4_1 BL BLB W_4_15_1 W_4_15_1_bar CIM_cell
X442 I415_inv O_4_15_2 WL_4_2 BL BLB W_4_15_2 W_4_15_2_bar CIM_cell
X443 I415_inv O_4_15_3 WL_4_3 BL BLB W_4_15_3 W_4_15_3_bar CIM_cell
X444 I415_inv O_4_15_4 WL_4_4 BL BLB W_4_15_4 W_4_15_4_bar CIM_cell
X445 I416_inv O_4_16_1 WL_4_1 BL BLB W_4_16_1 W_4_16_1_bar CIM_cell
X446 I416_inv O_4_16_2 WL_4_2 BL BLB W_4_16_2 W_4_16_2_bar CIM_cell
X447 I416_inv O_4_16_3 WL_4_3 BL BLB W_4_16_3 W_4_16_3_bar CIM_cell
X448 I416_inv O_4_16_4 WL_4_4 BL BLB W_4_16_4 W_4_16_4_bar CIM_cell
X449 I417_inv O_4_17_1 WL_4_1 BL BLB W_4_17_1 W_4_17_1_bar CIM_cell
X450 I417_inv O_4_17_2 WL_4_2 BL BLB W_4_17_2 W_4_17_2_bar CIM_cell
X451 I417_inv O_4_17_3 WL_4_3 BL BLB W_4_17_3 W_4_17_3_bar CIM_cell
X452 I417_inv O_4_17_4 WL_4_4 BL BLB W_4_17_4 W_4_17_4_bar CIM_cell
X453 I418_inv O_4_18_1 WL_4_1 BL BLB W_4_18_1 W_4_18_1_bar CIM_cell
X454 I418_inv O_4_18_2 WL_4_2 BL BLB W_4_18_2 W_4_18_2_bar CIM_cell
X455 I418_inv O_4_18_3 WL_4_3 BL BLB W_4_18_3 W_4_18_3_bar CIM_cell
X456 I418_inv O_4_18_4 WL_4_4 BL BLB W_4_18_4 W_4_18_4_bar CIM_cell
X457 I419_inv O_4_19_1 WL_4_1 BL BLB W_4_19_1 W_4_19_1_bar CIM_cell
X458 I419_inv O_4_19_2 WL_4_2 BL BLB W_4_19_2 W_4_19_2_bar CIM_cell
X459 I419_inv O_4_19_3 WL_4_3 BL BLB W_4_19_3 W_4_19_3_bar CIM_cell
X460 I419_inv O_4_19_4 WL_4_4 BL BLB W_4_19_4 W_4_19_4_bar CIM_cell
X461 I420_inv O_4_20_1 WL_4_1 BL BLB W_4_20_1 W_4_20_1_bar CIM_cell
X462 I420_inv O_4_20_2 WL_4_2 BL BLB W_4_20_2 W_4_20_2_bar CIM_cell
X463 I420_inv O_4_20_3 WL_4_3 BL BLB W_4_20_3 W_4_20_3_bar CIM_cell
X464 I420_inv O_4_20_4 WL_4_4 BL BLB W_4_20_4 W_4_20_4_bar CIM_cell
X465 I421_inv O_4_21_1 WL_4_1 BL BLB W_4_21_1 W_4_21_1_bar CIM_cell
X466 I421_inv O_4_21_2 WL_4_2 BL BLB W_4_21_2 W_4_21_2_bar CIM_cell
X467 I421_inv O_4_21_3 WL_4_3 BL BLB W_4_21_3 W_4_21_3_bar CIM_cell
X468 I421_inv O_4_21_4 WL_4_4 BL BLB W_4_21_4 W_4_21_4_bar CIM_cell
X469 I422_inv O_4_22_1 WL_4_1 BL BLB W_4_22_1 W_4_22_1_bar CIM_cell
X470 I422_inv O_4_22_2 WL_4_2 BL BLB W_4_22_2 W_4_22_2_bar CIM_cell
X471 I422_inv O_4_22_3 WL_4_3 BL BLB W_4_22_3 W_4_22_3_bar CIM_cell
X472 I422_inv O_4_22_4 WL_4_4 BL BLB W_4_22_4 W_4_22_4_bar CIM_cell
X473 I423_inv O_4_23_1 WL_4_1 BL BLB W_4_23_1 W_4_23_1_bar CIM_cell
X474 I423_inv O_4_23_2 WL_4_2 BL BLB W_4_23_2 W_4_23_2_bar CIM_cell
X475 I423_inv O_4_23_3 WL_4_3 BL BLB W_4_23_3 W_4_23_3_bar CIM_cell
X476 I423_inv O_4_23_4 WL_4_4 BL BLB W_4_23_4 W_4_23_4_bar CIM_cell
X477 I424_inv O_4_24_1 WL_4_1 BL BLB W_4_24_1 W_4_24_1_bar CIM_cell
X478 I424_inv O_4_24_2 WL_4_2 BL BLB W_4_24_2 W_4_24_2_bar CIM_cell
X479 I424_inv O_4_24_3 WL_4_3 BL BLB W_4_24_3 W_4_24_3_bar CIM_cell
X480 I424_inv O_4_24_4 WL_4_4 BL BLB W_4_24_4 W_4_24_4_bar CIM_cell
X481 I425_inv O_4_25_1 WL_4_1 BL BLB W_4_25_1 W_4_25_1_bar CIM_cell
X482 I425_inv O_4_25_2 WL_4_2 BL BLB W_4_25_2 W_4_25_2_bar CIM_cell
X483 I425_inv O_4_25_3 WL_4_3 BL BLB W_4_25_3 W_4_25_3_bar CIM_cell
X484 I425_inv O_4_25_4 WL_4_4 BL BLB W_4_25_4 W_4_25_4_bar CIM_cell
X485 I426_inv O_4_26_1 WL_4_1 BL BLB W_4_26_1 W_4_26_1_bar CIM_cell
X486 I426_inv O_4_26_2 WL_4_2 BL BLB W_4_26_2 W_4_26_2_bar CIM_cell
X487 I426_inv O_4_26_3 WL_4_3 BL BLB W_4_26_3 W_4_26_3_bar CIM_cell
X488 I426_inv O_4_26_4 WL_4_4 BL BLB W_4_26_4 W_4_26_4_bar CIM_cell
X489 I427_inv O_4_27_1 WL_4_1 BL BLB W_4_27_1 W_4_27_1_bar CIM_cell
X490 I427_inv O_4_27_2 WL_4_2 BL BLB W_4_27_2 W_4_27_2_bar CIM_cell
X491 I427_inv O_4_27_3 WL_4_3 BL BLB W_4_27_3 W_4_27_3_bar CIM_cell
X492 I427_inv O_4_27_4 WL_4_4 BL BLB W_4_27_4 W_4_27_4_bar CIM_cell
X493 I428_inv O_4_28_1 WL_4_1 BL BLB W_4_28_1 W_4_28_1_bar CIM_cell
X494 I428_inv O_4_28_2 WL_4_2 BL BLB W_4_28_2 W_4_28_2_bar CIM_cell
X495 I428_inv O_4_28_3 WL_4_3 BL BLB W_4_28_3 W_4_28_3_bar CIM_cell
X496 I428_inv O_4_28_4 WL_4_4 BL BLB W_4_28_4 W_4_28_4_bar CIM_cell
X497 I429_inv O_4_29_1 WL_4_1 BL BLB W_4_29_1 W_4_29_1_bar CIM_cell
X498 I429_inv O_4_29_2 WL_4_2 BL BLB W_4_29_2 W_4_29_2_bar CIM_cell
X499 I429_inv O_4_29_3 WL_4_3 BL BLB W_4_29_3 W_4_29_3_bar CIM_cell
X500 I429_inv O_4_29_4 WL_4_4 BL BLB W_4_29_4 W_4_29_4_bar CIM_cell
X501 I430_inv O_4_30_1 WL_4_1 BL BLB W_4_30_1 W_4_30_1_bar CIM_cell
X502 I430_inv O_4_30_2 WL_4_2 BL BLB W_4_30_2 W_4_30_2_bar CIM_cell
X503 I430_inv O_4_30_3 WL_4_3 BL BLB W_4_30_3 W_4_30_3_bar CIM_cell
X504 I430_inv O_4_30_4 WL_4_4 BL BLB W_4_30_4 W_4_30_4_bar CIM_cell
X505 I431_inv O_4_31_1 WL_4_1 BL BLB W_4_31_1 W_4_31_1_bar CIM_cell
X506 I431_inv O_4_31_2 WL_4_2 BL BLB W_4_31_2 W_4_31_2_bar CIM_cell
X507 I431_inv O_4_31_3 WL_4_3 BL BLB W_4_31_3 W_4_31_3_bar CIM_cell
X508 I431_inv O_4_31_4 WL_4_4 BL BLB W_4_31_4 W_4_31_4_bar CIM_cell
X509 I432_inv O_4_32_1 WL_4_1 BL BLB W_4_32_1 W_4_32_1_bar CIM_cell
X510 I432_inv O_4_32_2 WL_4_2 BL BLB W_4_32_2 W_4_32_2_bar CIM_cell
X511 I432_inv O_4_32_3 WL_4_3 BL BLB W_4_32_3 W_4_32_3_bar CIM_cell
X512 I432_inv O_4_32_4 WL_4_4 BL BLB W_4_32_4 W_4_32_4_bar CIM_cell


X513 GND VDD O_1_1_4 O_1_1_3 O_1_1_2 O_1_1_1 O_1_2_4 O_1_2_3 O_1_2_2 O_1_2_1 O_1_3_4 O_1_3_3 O_1_3_2 O_1_3_1 O_1_4_4 O_1_4_3 O_1_4_2 O_1_4_1 
+ O_1_5_4 O_1_5_3 O_1_5_2 O_1_5_1 O_1_6_4 O_1_6_3 O_1_6_2 O_1_6_1 O_1_7_4 O_1_7_3 O_1_7_2 O_1_7_1 O_1_8_4 O_1_8_3 O_1_8_2 O_1_8_1
+ O_1_9_4 O_1_9_3 O_1_9_2 O_1_9_1 O_1_10_4 O_1_10_3 O_1_10_2 O_1_10_1 O_1_11_4 O_1_11_3 O_1_11_2 O_1_11_1 O_1_12_4 O_1_12_3 O_1_12_2 O_1_12_1 
+ O_1_13_4 O_1_13_3 O_1_13_2 O_1_13_1 O_1_14_4 O_1_14_3 O_1_14_2 O_1_14_1 O_1_15_4 O_1_15_3 O_1_15_2 O_1_15_1 O_1_16_4 O_1_16_3 O_1_16_2 O_1_16_1 
+ O_1_17_4 O_1_17_3 O_1_17_2 O_1_17_1 O_1_18_4 O_1_18_3 O_1_18_2 O_1_18_1 O_1_19_4 O_1_19_3 O_1_19_2 O_1_19_1 O_1_20_4 O_1_20_3 O_1_20_2 O_1_20_1 
+ O_1_21_4 O_1_21_3 O_1_21_2 O_1_21_1 O_1_22_4 O_1_22_3 O_1_22_2 O_1_22_1 O_1_23_4 O_1_23_3 O_1_23_2 O_1_23_1 O_1_24_4 O_1_24_3 O_1_24_2 O_1_24_1 
+ O_1_25_4 O_1_25_3 O_1_25_2 O_1_25_1 O_1_26_4 O_1_26_3 O_1_26_2 O_1_26_1 O_1_27_4 O_1_27_3 O_1_27_2 O_1_27_1 O_1_28_4 O_1_28_3 O_1_28_2 O_1_28_1 
+ O_1_29_4 O_1_29_3 O_1_29_2 O_1_29_1 O_1_30_4 O_1_30_3 O_1_30_2 O_1_30_1 O_1_31_4 O_1_31_3 O_1_31_2 O_1_31_1 O_1_32_4 O_1_32_3 O_1_32_2 O_1_32_1 
​+ partial_sum_12_1 partial_sum_11_1 partial_sum_10_1 partial_sum_9_1 partial_sum_8_1 partial_sum_7_1 partial_sum_6_1 partial_sum_5_1 partial_sum_4_1 partial_sum_3_1 partial_sum_2_1 partial_sum_1_1 partial_sum_0_1 Adder_tree

X514 GND VDD O_2_1_4 O_2_1_3 O_2_1_2 O_2_1_1 O_2_2_4 O_2_2_3 O_2_2_2 O_2_2_1 O_2_3_4 O_2_3_3 O_2_3_2 O_2_3_1 O_2_4_4 O_2_4_3 O_2_4_2 O_2_4_1 
+ O_2_5_4 O_2_5_3 O_2_5_2 O_2_5_1 O_2_6_4 O_2_6_3 O_2_6_2 O_2_6_1 O_2_7_4 O_2_7_3 O_2_7_2 O_2_7_1 O_2_8_4 O_2_8_3 O_2_8_2 O_2_8_1 
+ O_2_9_4 O_2_9_3 O_2_9_2 O_2_9_1 O_2_10_4 O_2_10_3 O_2_10_2 O_2_10_1 O_2_11_4 O_2_11_3 O_2_11_2 O_2_11_1 O_2_12_4 O_2_12_3 O_2_12_2 O_2_12_1 
+ O_2_13_4 O_2_13_3 O_2_13_2 O_2_13_1 O_2_14_4 O_2_14_3 O_2_14_2 O_2_14_1 O_2_15_4 O_2_15_3 O_2_15_2 O_2_15_1 O_2_16_4 O_2_16_3 O_2_16_2 O_2_16_1 
+ O_2_17_4 O_2_17_3 O_2_17_2 O_2_17_1 O_2_18_4 O_2_18_3 O_2_18_2 O_2_18_1 O_2_19_4 O_2_19_3 O_2_19_2 O_2_19_1 O_2_20_4 O_2_20_3 O_2_20_2 O_2_20_1
+ O_2_21_4 O_2_21_3 O_2_21_2 O_2_21_1 O_2_22_4 O_2_22_3 O_2_22_2 O_2_22_1 O_2_23_4 O_2_23_3 O_2_23_2 O_2_23_1 O_2_24_4 O_2_24_3 O_2_24_2 O_2_24_1 
+ O_2_25_4 O_2_25_3 O_2_25_2 O_2_25_1 O_2_26_4 O_2_26_3 O_2_26_2 O_2_26_1 O_2_27_4 O_2_27_3 O_2_27_2 O_2_27_1 O_2_28_4 O_2_28_3 O_2_28_2 O_2_28_1 
+ O_2_29_4 O_2_29_3 O_2_29_2 O_2_29_1 O_2_30_4 O_2_30_3 O_2_30_2 O_2_30_1 O_2_31_4 O_2_31_3 O_2_31_2 O_2_31_1 O_2_32_4 O_2_32_3 O_2_32_2 O_2_32_1 
+ partial_sum_12_2 partial_sum_11_2 partial_sum_10_2 partial_sum_9_2 partial_sum_8_2 partial_sum_7_2 partial_sum_6_2 partial_sum_5_2 partial_sum_4_2 partial_sum_3_2 partial_sum_2_2 partial_sum_1_2 partial_sum_0_2 Adder_tree

X515 GND VDD O_3_1_4 O_3_1_3 O_3_1_2 O_3_1_1 O_3_2_4 O_3_2_3 O_3_2_2 O_3_2_1 O_3_3_4 O_3_3_3 O_3_3_2 O_3_3_1 O_3_4_4 O_3_4_3 O_3_4_2 O_3_4_1 
+ O_3_5_4 O_3_5_3 O_3_5_2 O_3_5_1 O_3_6_4 O_3_6_3 O_3_6_2 O_3_6_1 O_3_7_4 O_3_7_3 O_3_7_2 O_3_7_1 O_3_8_4 O_3_8_3 O_3_8_2 O_3_8_1 
+ O_3_9_4 O_3_9_3 O_3_9_2 O_3_9_1 O_3_10_4 O_3_10_3 O_3_10_2 O_3_10_1 O_3_11_4 O_3_11_3 O_3_11_2 O_3_11_1 O_3_12_4 O_3_12_3 O_3_12_2 O_3_12_1 
+ O_3_13_4 O_3_13_3 O_3_13_2 O_3_13_1 O_3_14_4 O_3_14_3 O_3_14_2 O_3_14_1 O_3_15_4 O_3_15_3 O_3_15_2 O_3_15_1 O_3_16_4 O_3_16_3 O_3_16_2 O_3_16_1 
+ O_3_17_4 O_3_17_3 O_3_17_2 O_3_17_1 O_3_18_4 O_3_18_3 O_3_18_2 O_3_18_1 O_3_19_4 O_3_19_3 O_3_19_2 O_3_19_1 O_3_20_4 O_3_20_3 O_3_20_2 O_3_20_1 
+ O_3_21_4 O_3_21_3 O_3_21_2 O_3_21_1 O_3_22_4 O_3_22_3 O_3_22_2 O_3_22_1 O_3_23_4 O_3_23_3 O_3_23_2 O_3_23_1 O_3_24_4 O_3_24_3 O_3_24_2 O_3_24_1 
+ O_3_25_4 O_3_25_3 O_3_25_2 O_3_25_1 O_3_26_4 O_3_26_3 O_3_26_2 O_3_26_1 O_3_27_4 O_3_27_3 O_3_27_2 O_3_27_1 O_3_28_4 O_3_28_3 O_3_28_2 O_3_28_1 
+ O_3_29_4 O_3_29_3 O_3_29_2 O_3_29_1 O_3_30_4 O_3_30_3 O_3_30_2 O_3_30_1 O_3_31_4 O_3_31_3 O_3_31_2 O_3_31_1 O_3_32_4 O_3_32_3 O_3_32_2 O_3_32_1 
+ partial_sum_12_3 partial_sum_11_3 partial_sum_10_3 partial_sum_9_3 partial_sum_8_3 partial_sum_7_3 partial_sum_6_3 partial_sum_5_3 partial_sum_4_3 partial_sum_3_3 partial_sum_2_3 partial_sum_1_3 partial_sum_0_3 Adder_tree

X516 GND VDD O_4_1_4 O_4_1_3 O_4_1_2 O_4_1_1 O_4_2_4 O_4_2_3 O_4_2_2 O_4_2_1 O_4_3_4 O_4_3_3 O_4_3_2 O_4_3_1 O_4_4_4 O_4_4_3 O_4_4_2 O_4_4_1 
+ O_4_5_4 O_4_5_3 O_4_5_2 O_4_5_1 O_4_6_4 O_4_6_3 O_4_6_2 O_4_6_1 O_4_7_4 O_4_7_3 O_4_7_2 O_4_7_1 O_4_8_4 O_4_8_3 O_4_8_2 O_4_8_1 
+ O_4_9_4 O_4_9_3 O_4_9_2 O_4_9_1 O_4_10_4 O_4_10_3 O_4_10_2 O_4_10_1 O_4_11_4 O_4_11_3 O_4_11_2 O_4_11_1 O_4_12_4 O_4_12_3 O_4_12_2 O_4_12_1 
+ O_4_13_4 O_4_13_3 O_4_13_2 O_4_13_1 O_4_14_4 O_4_14_3 O_4_14_2 O_4_14_1 O_4_15_4 O_4_15_3 O_4_15_2 O_4_15_1 O_4_16_4 O_4_16_3 O_4_16_2 O_4_16_1 
+ O_4_17_4 O_4_17_3 O_4_17_2 O_4_17_1 O_4_18_4 O_4_18_3 O_4_18_2 O_4_18_1 O_4_19_4 O_4_19_3 O_4_19_2 O_4_19_1 O_4_20_4 O_4_20_3 O_4_20_2 O_4_20_1 
+ O_4_21_4 O_4_21_3 O_4_21_2 O_4_21_1 O_4_22_4 O_4_22_3 O_4_22_2 O_4_22_1 O_4_23_4 O_4_23_3 O_4_23_2 O_4_23_1 O_4_24_4 O_4_24_3 O_4_24_2 O_4_24_1 
+ O_4_25_4 O_4_25_3 O_4_25_2 O_4_25_1 O_4_26_4 O_4_26_3 O_4_26_2 O_4_26_1 O_4_27_4 O_4_27_3 O_4_27_2 O_4_27_1 O_4_28_4 O_4_28_3 O_4_28_2 O_4_28_1 
+ O_4_29_4 O_4_29_3 O_4_29_2 O_4_29_1 O_4_30_4 O_4_30_3 O_4_30_2 O_4_30_1 O_4_31_4 O_4_31_3 O_4_31_2 O_4_31_1 O_4_32_4 O_4_32_3 O_4_32_2 O_4_32_1 
+ partial_sum_12_4 partial_sum_11_4 partial_sum_10_4 partial_sum_9_4 partial_sum_8_4 partial_sum_7_4 partial_sum_6_4 partial_sum_5_4 partial_sum_4_4 partial_sum_3_4 partial_sum_2_4 partial_sum_1_4 partial_sum_0_4 Adder_tree


X517 GND VDD clk rst_n in_valid partial_sum_12_1 partial_sum_11_1 partial_sum_10_1 partial_sum_9_1 partial_sum_8_1 partial_sum_7_1 partial_sum_6_1 partial_sum_5_1 partial_sum_4_1 partial_sum_3_1 partial_sum_2_1 partial_sum_1_1 partial_sum_0_1 Out_1[12]  Out_1[11]  Out_1[10]  Out_1[9]  Out_1[8]  Out_1[7]  Out_1[6]  Out_1[5]  Out_1[4]  Out_1[3]  Out_1[2]  Out_1[1]  Out_1[0]  Accumulator          
*X518 GND VDD clk rst_n in_valid partial_sum_12_2 partial_sum_11_2 partial_sum_10_2 partial_sum_9_2 partial_sum_8_2 partial_sum_7_2 partial_sum_6_2 partial_sum_5_2 partial_sum_4_2 partial_sum_3_2 partial_sum_2_2 partial_sum_1_2 partial_sum_0_2  Output_12_2 Output_11_2 Output_10_2 Output_9_2 Output_8_2 Output_7_2 Output_6_2 Output_5_2 Output_4_2 Output_3_2 Output_2_2 Output_1_2 Output_0_2  Accumulator 
*X519 GND VDD clk rst_n in_valid partial_sum_12_3 partial_sum_11_3 partial_sum_10_3 partial_sum_9_3 partial_sum_8_3 partial_sum_7_3 partial_sum_6_3 partial_sum_5_3 partial_sum_4_3 partial_sum_3_3 partial_sum_2_3 partial_sum_1_3 partial_sum_0_3  Output_12_3 Output_11_3 Output_10_3 Output_9_3 Output_8_3 Output_7_3 Output_6_3 Output_5_3 Output_4_3 Output_3_3 Output_2_3 Output_1_3 Output_0_3  Accumulator 
*X520 GND VDD clk rst_n in_valid partial_sum_12_4 partial_sum_11_4 partial_sum_10_4 partial_sum_9_4 partial_sum_8_4 partial_sum_7_4 partial_sum_6_4 partial_sum_5_4 partial_sum_4_4 partial_sum_3_4 partial_sum_2_4 partial_sum_1_4 partial_sum_0_4  Output_12_4 Output_11_4 Output_10_4 Output_9_4 Output_8_4 Output_7_4 Output_6_4 Output_5_4 Output_4_4 Output_3_4 Output_2_4 Output_1_4 Output_0_4  Accumulator 

***-----------------------***
***      sub-circuit      ***
***-----------------------***

* // QB : weight 
* // input 
* // output 
* .subckt CIM_cell Input Output WL BL BLB q qb
*     X01 WL BL BLB q qb SRAM_6T
*     X02 qb Input Output NOR_2
* .ends

.subckt CIM_cell Input Output WL BL BLB q qb
    X01 WL BL BLB q qb SRAM_6T
    X02 qb Input Output NOR_2
.ends


.subckt SRAM_6T WL BL BLB q qb
    MP1 q   qb  VDD VDD pmos_sram m=1
    MP2 qb  q   VDD VDD pmos_sram m=1
    MN1 q   qb  GND GND nmos_sram m=1
    MN2 qb  q   GND GND nmos_sram m=1
    MN3 BL  WL  q   GND nmos_sram m=1
    MN4 qb  WL  BLB GND nmos_sram m=1
.ends

.subckt NOR_2 A B Y
    MP1 N1  A   VDD VDD pmos_lvt m=1
    MP2 Y   B   N1  VDD pmos_lvt m=1
    MN1 Y   A   GND GND nmos_lvt m=1
    MN2 Y   B   GND GND nmos_lvt m=1
.ends

.subckt Buffer in out
    X_INV1 in   in_b INV
    X_INV2 in_b out  INV
.ends

.subckt INV in out
    Mp  out  in  VDD  VDD  pmos_lvt  m=1
    Mn  out  in  GND  GND  nmos_lvt  m=1
.ends

* Example .IC file for initializing SRAM weights
.IC V(W_1_1_1) = 1 V(W_1_1_1_bar) = 0
.IC V(W_1_1_2) = 1 V(W_1_1_2_bar) = 0
.IC V(W_1_1_3) = 1 V(W_1_1_3_bar) = 0
.IC V(W_1_1_4) = 1 V(W_1_1_4_bar) = 0
.IC V(W_1_2_1) = 1 V(W_1_2_1_bar) = 0
.IC V(W_1_2_2) = 1 V(W_1_2_2_bar) = 0
.IC V(W_1_2_3) = 1 V(W_1_2_3_bar) = 0
.IC V(W_1_2_4) = 1 V(W_1_2_4_bar) = 0
.IC V(W_1_3_1) = 0 V(W_1_3_1_bar) = 1
.IC V(W_1_3_2) = 0 V(W_1_3_2_bar) = 1
.IC V(W_1_3_3) = 0 V(W_1_3_3_bar) = 1
.IC V(W_1_3_4) = 0 V(W_1_3_4_bar) = 1
.IC V(W_1_4_1) = 0 V(W_1_4_1_bar) = 1
.IC V(W_1_4_2) = 1 V(W_1_4_2_bar) = 0
.IC V(W_1_4_3) = 0 V(W_1_4_3_bar) = 1
.IC V(W_1_4_4) = 1 V(W_1_4_4_bar) = 0
.IC V(W_1_5_1) = 0 V(W_1_5_1_bar) = 1
.IC V(W_1_5_2) = 0 V(W_1_5_2_bar) = 1
.IC V(W_1_5_3) = 1 V(W_1_5_3_bar) = 0
.IC V(W_1_5_4) = 0 V(W_1_5_4_bar) = 1
.IC V(W_1_6_1) = 0 V(W_1_6_1_bar) = 1
.IC V(W_1_6_2) = 0 V(W_1_6_2_bar) = 1
.IC V(W_1_6_3) = 1 V(W_1_6_3_bar) = 0
.IC V(W_1_6_4) = 0 V(W_1_6_4_bar) = 1
.IC V(W_1_7_1) = 0 V(W_1_7_1_bar) = 1
.IC V(W_1_7_2) = 1 V(W_1_7_2_bar) = 0
.IC V(W_1_7_3) = 1 V(W_1_7_3_bar) = 0
.IC V(W_1_7_4) = 1 V(W_1_7_4_bar) = 0
.IC V(W_1_8_1) = 1 V(W_1_8_1_bar) = 0
.IC V(W_1_8_2) = 1 V(W_1_8_2_bar) = 0
.IC V(W_1_8_3) = 0 V(W_1_8_3_bar) = 1
.IC V(W_1_8_4) = 0 V(W_1_8_4_bar) = 1
.IC V(W_1_9_1) = 1 V(W_1_9_1_bar) = 0
.IC V(W_1_9_2) = 1 V(W_1_9_2_bar) = 0
.IC V(W_1_9_3) = 0 V(W_1_9_3_bar) = 1
.IC V(W_1_9_4) = 1 V(W_1_9_4_bar) = 0
.IC V(W_1_10_1) = 1 V(W_1_10_1_bar) = 0
.IC V(W_1_10_2) = 0 V(W_1_10_2_bar) = 1
.IC V(W_1_10_3) = 0 V(W_1_10_3_bar) = 1
.IC V(W_1_10_4) = 1 V(W_1_10_4_bar) = 0
.IC V(W_1_11_1) = 1 V(W_1_11_1_bar) = 0
.IC V(W_1_11_2) = 1 V(W_1_11_2_bar) = 0
.IC V(W_1_11_3) = 0 V(W_1_11_3_bar) = 1
.IC V(W_1_11_4) = 1 V(W_1_11_4_bar) = 0
.IC V(W_1_12_1) = 1 V(W_1_12_1_bar) = 0
.IC V(W_1_12_2) = 1 V(W_1_12_2_bar) = 0
.IC V(W_1_12_3) = 1 V(W_1_12_3_bar) = 0
.IC V(W_1_12_4) = 1 V(W_1_12_4_bar) = 0
.IC V(W_1_13_1) = 1 V(W_1_13_1_bar) = 0
.IC V(W_1_13_2) = 0 V(W_1_13_2_bar) = 1
.IC V(W_1_13_3) = 0 V(W_1_13_3_bar) = 1
.IC V(W_1_13_4) = 0 V(W_1_13_4_bar) = 1
.IC V(W_1_14_1) = 1 V(W_1_14_1_bar) = 0
.IC V(W_1_14_2) = 0 V(W_1_14_2_bar) = 1
.IC V(W_1_14_3) = 0 V(W_1_14_3_bar) = 1
.IC V(W_1_14_4) = 1 V(W_1_14_4_bar) = 0
.IC V(W_1_15_1) = 0 V(W_1_15_1_bar) = 1
.IC V(W_1_15_2) = 0 V(W_1_15_2_bar) = 1
.IC V(W_1_15_3) = 0 V(W_1_15_3_bar) = 1
.IC V(W_1_15_4) = 0 V(W_1_15_4_bar) = 1
.IC V(W_1_16_1) = 1 V(W_1_16_1_bar) = 0
.IC V(W_1_16_2) = 0 V(W_1_16_2_bar) = 1
.IC V(W_1_16_3) = 0 V(W_1_16_3_bar) = 1
.IC V(W_1_16_4) = 0 V(W_1_16_4_bar) = 1
.IC V(W_1_17_1) = 1 V(W_1_17_1_bar) = 0
.IC V(W_1_17_2) = 0 V(W_1_17_2_bar) = 1
.IC V(W_1_17_3) = 0 V(W_1_17_3_bar) = 1
.IC V(W_1_17_4) = 1 V(W_1_17_4_bar) = 0
.IC V(W_1_18_1) = 1 V(W_1_18_1_bar) = 0
.IC V(W_1_18_2) = 1 V(W_1_18_2_bar) = 0
.IC V(W_1_18_3) = 1 V(W_1_18_3_bar) = 0
.IC V(W_1_18_4) = 0 V(W_1_18_4_bar) = 1
.IC V(W_1_19_1) = 1 V(W_1_19_1_bar) = 0
.IC V(W_1_19_2) = 1 V(W_1_19_2_bar) = 0
.IC V(W_1_19_3) = 1 V(W_1_19_3_bar) = 0
.IC V(W_1_19_4) = 1 V(W_1_19_4_bar) = 0
.IC V(W_1_20_1) = 0 V(W_1_20_1_bar) = 1
.IC V(W_1_20_2) = 0 V(W_1_20_2_bar) = 1
.IC V(W_1_20_3) = 1 V(W_1_20_3_bar) = 0
.IC V(W_1_20_4) = 0 V(W_1_20_4_bar) = 1
.IC V(W_1_21_1) = 1 V(W_1_21_1_bar) = 0
.IC V(W_1_21_2) = 1 V(W_1_21_2_bar) = 0
.IC V(W_1_21_3) = 1 V(W_1_21_3_bar) = 0
.IC V(W_1_21_4) = 1 V(W_1_21_4_bar) = 0
.IC V(W_1_22_1) = 0 V(W_1_22_1_bar) = 1
.IC V(W_1_22_2) = 1 V(W_1_22_2_bar) = 0
.IC V(W_1_22_3) = 1 V(W_1_22_3_bar) = 0
.IC V(W_1_22_4) = 0 V(W_1_22_4_bar) = 1
.IC V(W_1_23_1) = 1 V(W_1_23_1_bar) = 0
.IC V(W_1_23_2) = 0 V(W_1_23_2_bar) = 1
.IC V(W_1_23_3) = 1 V(W_1_23_3_bar) = 0
.IC V(W_1_23_4) = 1 V(W_1_23_4_bar) = 0
.IC V(W_1_24_1) = 0 V(W_1_24_1_bar) = 1
.IC V(W_1_24_2) = 1 V(W_1_24_2_bar) = 0
.IC V(W_1_24_3) = 0 V(W_1_24_3_bar) = 1
.IC V(W_1_24_4) = 1 V(W_1_24_4_bar) = 0
.IC V(W_1_25_1) = 1 V(W_1_25_1_bar) = 0
.IC V(W_1_25_2) = 1 V(W_1_25_2_bar) = 0
.IC V(W_1_25_3) = 1 V(W_1_25_3_bar) = 0
.IC V(W_1_25_4) = 1 V(W_1_25_4_bar) = 0
.IC V(W_1_26_1) = 1 V(W_1_26_1_bar) = 0
.IC V(W_1_26_2) = 0 V(W_1_26_2_bar) = 1
.IC V(W_1_26_3) = 1 V(W_1_26_3_bar) = 0
.IC V(W_1_26_4) = 0 V(W_1_26_4_bar) = 1
.IC V(W_1_27_1) = 1 V(W_1_27_1_bar) = 0
.IC V(W_1_27_2) = 1 V(W_1_27_2_bar) = 0
.IC V(W_1_27_3) = 1 V(W_1_27_3_bar) = 0
.IC V(W_1_27_4) = 0 V(W_1_27_4_bar) = 1
.IC V(W_1_28_1) = 0 V(W_1_28_1_bar) = 1
.IC V(W_1_28_2) = 0 V(W_1_28_2_bar) = 1
.IC V(W_1_28_3) = 1 V(W_1_28_3_bar) = 0
.IC V(W_1_28_4) = 1 V(W_1_28_4_bar) = 0
.IC V(W_1_29_1) = 0 V(W_1_29_1_bar) = 1
.IC V(W_1_29_2) = 1 V(W_1_29_2_bar) = 0
.IC V(W_1_29_3) = 1 V(W_1_29_3_bar) = 0
.IC V(W_1_29_4) = 0 V(W_1_29_4_bar) = 1
.IC V(W_1_30_1) = 0 V(W_1_30_1_bar) = 1
.IC V(W_1_30_2) = 0 V(W_1_30_2_bar) = 1
.IC V(W_1_30_3) = 1 V(W_1_30_3_bar) = 0
.IC V(W_1_30_4) = 0 V(W_1_30_4_bar) = 1
.IC V(W_1_31_1) = 1 V(W_1_31_1_bar) = 0
.IC V(W_1_31_2) = 1 V(W_1_31_2_bar) = 0
.IC V(W_1_31_3) = 1 V(W_1_31_3_bar) = 0
.IC V(W_1_31_4) = 0 V(W_1_31_4_bar) = 1
.IC V(W_1_32_1) = 0 V(W_1_32_1_bar) = 1
.IC V(W_1_32_2) = 1 V(W_1_32_2_bar) = 0
.IC V(W_1_32_3) = 1 V(W_1_32_3_bar) = 0
.IC V(W_1_32_4) = 1 V(W_1_32_4_bar) = 0
.IC V(W_2_1_1) = 1 V(W_2_1_1_bar) = 0
.IC V(W_2_1_2) = 0 V(W_2_1_2_bar) = 1
.IC V(W_2_1_3) = 1 V(W_2_1_3_bar) = 0
.IC V(W_2_1_4) = 1 V(W_2_1_4_bar) = 0
.IC V(W_2_2_1) = 1 V(W_2_2_1_bar) = 0
.IC V(W_2_2_2) = 0 V(W_2_2_2_bar) = 1
.IC V(W_2_2_3) = 0 V(W_2_2_3_bar) = 1
.IC V(W_2_2_4) = 0 V(W_2_2_4_bar) = 1
.IC V(W_2_3_1) = 0 V(W_2_3_1_bar) = 1
.IC V(W_2_3_2) = 0 V(W_2_3_2_bar) = 1
.IC V(W_2_3_3) = 1 V(W_2_3_3_bar) = 0
.IC V(W_2_3_4) = 0 V(W_2_3_4_bar) = 1
.IC V(W_2_4_1) = 0 V(W_2_4_1_bar) = 1
.IC V(W_2_4_2) = 0 V(W_2_4_2_bar) = 1
.IC V(W_2_4_3) = 0 V(W_2_4_3_bar) = 1
.IC V(W_2_4_4) = 1 V(W_2_4_4_bar) = 0
.IC V(W_2_5_1) = 0 V(W_2_5_1_bar) = 1
.IC V(W_2_5_2) = 1 V(W_2_5_2_bar) = 0
.IC V(W_2_5_3) = 0 V(W_2_5_3_bar) = 1
.IC V(W_2_5_4) = 1 V(W_2_5_4_bar) = 0
.IC V(W_2_6_1) = 0 V(W_2_6_1_bar) = 1
.IC V(W_2_6_2) = 0 V(W_2_6_2_bar) = 1
.IC V(W_2_6_3) = 0 V(W_2_6_3_bar) = 1
.IC V(W_2_6_4) = 1 V(W_2_6_4_bar) = 0
.IC V(W_2_7_1) = 1 V(W_2_7_1_bar) = 0
.IC V(W_2_7_2) = 0 V(W_2_7_2_bar) = 1
.IC V(W_2_7_3) = 0 V(W_2_7_3_bar) = 1
.IC V(W_2_7_4) = 0 V(W_2_7_4_bar) = 1
.IC V(W_2_8_1) = 1 V(W_2_8_1_bar) = 0
.IC V(W_2_8_2) = 0 V(W_2_8_2_bar) = 1
.IC V(W_2_8_3) = 0 V(W_2_8_3_bar) = 1
.IC V(W_2_8_4) = 1 V(W_2_8_4_bar) = 0
.IC V(W_2_9_1) = 0 V(W_2_9_1_bar) = 1
.IC V(W_2_9_2) = 1 V(W_2_9_2_bar) = 0
.IC V(W_2_9_3) = 0 V(W_2_9_3_bar) = 1
.IC V(W_2_9_4) = 1 V(W_2_9_4_bar) = 0
.IC V(W_2_10_1) = 0 V(W_2_10_1_bar) = 1
.IC V(W_2_10_2) = 0 V(W_2_10_2_bar) = 1
.IC V(W_2_10_3) = 0 V(W_2_10_3_bar) = 1
.IC V(W_2_10_4) = 0 V(W_2_10_4_bar) = 1
.IC V(W_2_11_1) = 0 V(W_2_11_1_bar) = 1
.IC V(W_2_11_2) = 0 V(W_2_11_2_bar) = 1
.IC V(W_2_11_3) = 1 V(W_2_11_3_bar) = 0
.IC V(W_2_11_4) = 0 V(W_2_11_4_bar) = 1
.IC V(W_2_12_1) = 0 V(W_2_12_1_bar) = 1
.IC V(W_2_12_2) = 0 V(W_2_12_2_bar) = 1
.IC V(W_2_12_3) = 0 V(W_2_12_3_bar) = 1
.IC V(W_2_12_4) = 0 V(W_2_12_4_bar) = 1
.IC V(W_2_13_1) = 0 V(W_2_13_1_bar) = 1
.IC V(W_2_13_2) = 0 V(W_2_13_2_bar) = 1
.IC V(W_2_13_3) = 1 V(W_2_13_3_bar) = 0
.IC V(W_2_13_4) = 1 V(W_2_13_4_bar) = 0
.IC V(W_2_14_1) = 0 V(W_2_14_1_bar) = 1
.IC V(W_2_14_2) = 0 V(W_2_14_2_bar) = 1
.IC V(W_2_14_3) = 1 V(W_2_14_3_bar) = 0
.IC V(W_2_14_4) = 0 V(W_2_14_4_bar) = 1
.IC V(W_2_15_1) = 0 V(W_2_15_1_bar) = 1
.IC V(W_2_15_2) = 0 V(W_2_15_2_bar) = 1
.IC V(W_2_15_3) = 1 V(W_2_15_3_bar) = 0
.IC V(W_2_15_4) = 1 V(W_2_15_4_bar) = 0
.IC V(W_2_16_1) = 0 V(W_2_16_1_bar) = 1
.IC V(W_2_16_2) = 1 V(W_2_16_2_bar) = 0
.IC V(W_2_16_3) = 0 V(W_2_16_3_bar) = 1
.IC V(W_2_16_4) = 1 V(W_2_16_4_bar) = 0
.IC V(W_2_17_1) = 0 V(W_2_17_1_bar) = 1
.IC V(W_2_17_2) = 1 V(W_2_17_2_bar) = 0
.IC V(W_2_17_3) = 1 V(W_2_17_3_bar) = 0
.IC V(W_2_17_4) = 0 V(W_2_17_4_bar) = 1
.IC V(W_2_18_1) = 0 V(W_2_18_1_bar) = 1
.IC V(W_2_18_2) = 1 V(W_2_18_2_bar) = 0
.IC V(W_2_18_3) = 0 V(W_2_18_3_bar) = 1
.IC V(W_2_18_4) = 0 V(W_2_18_4_bar) = 1
.IC V(W_2_19_1) = 1 V(W_2_19_1_bar) = 0
.IC V(W_2_19_2) = 1 V(W_2_19_2_bar) = 0
.IC V(W_2_19_3) = 0 V(W_2_19_3_bar) = 1
.IC V(W_2_19_4) = 1 V(W_2_19_4_bar) = 0
.IC V(W_2_20_1) = 1 V(W_2_20_1_bar) = 0
.IC V(W_2_20_2) = 1 V(W_2_20_2_bar) = 0
.IC V(W_2_20_3) = 0 V(W_2_20_3_bar) = 1
.IC V(W_2_20_4) = 1 V(W_2_20_4_bar) = 0
.IC V(W_2_21_1) = 0 V(W_2_21_1_bar) = 1
.IC V(W_2_21_2) = 1 V(W_2_21_2_bar) = 0
.IC V(W_2_21_3) = 0 V(W_2_21_3_bar) = 1
.IC V(W_2_21_4) = 1 V(W_2_21_4_bar) = 0
.IC V(W_2_22_1) = 0 V(W_2_22_1_bar) = 1
.IC V(W_2_22_2) = 0 V(W_2_22_2_bar) = 1
.IC V(W_2_22_3) = 0 V(W_2_22_3_bar) = 1
.IC V(W_2_22_4) = 0 V(W_2_22_4_bar) = 1
.IC V(W_2_23_1) = 0 V(W_2_23_1_bar) = 1
.IC V(W_2_23_2) = 1 V(W_2_23_2_bar) = 0
.IC V(W_2_23_3) = 1 V(W_2_23_3_bar) = 0
.IC V(W_2_23_4) = 0 V(W_2_23_4_bar) = 1
.IC V(W_2_24_1) = 0 V(W_2_24_1_bar) = 1
.IC V(W_2_24_2) = 0 V(W_2_24_2_bar) = 1
.IC V(W_2_24_3) = 1 V(W_2_24_3_bar) = 0
.IC V(W_2_24_4) = 1 V(W_2_24_4_bar) = 0
.IC V(W_2_25_1) = 1 V(W_2_25_1_bar) = 0
.IC V(W_2_25_2) = 0 V(W_2_25_2_bar) = 1
.IC V(W_2_25_3) = 0 V(W_2_25_3_bar) = 1
.IC V(W_2_25_4) = 0 V(W_2_25_4_bar) = 1
.IC V(W_2_26_1) = 1 V(W_2_26_1_bar) = 0
.IC V(W_2_26_2) = 0 V(W_2_26_2_bar) = 1
.IC V(W_2_26_3) = 1 V(W_2_26_3_bar) = 0
.IC V(W_2_26_4) = 1 V(W_2_26_4_bar) = 0
.IC V(W_2_27_1) = 1 V(W_2_27_1_bar) = 0
.IC V(W_2_27_2) = 1 V(W_2_27_2_bar) = 0
.IC V(W_2_27_3) = 0 V(W_2_27_3_bar) = 1
.IC V(W_2_27_4) = 1 V(W_2_27_4_bar) = 0
.IC V(W_2_28_1) = 0 V(W_2_28_1_bar) = 1
.IC V(W_2_28_2) = 0 V(W_2_28_2_bar) = 1
.IC V(W_2_28_3) = 0 V(W_2_28_3_bar) = 1
.IC V(W_2_28_4) = 1 V(W_2_28_4_bar) = 0
.IC V(W_2_29_1) = 0 V(W_2_29_1_bar) = 1
.IC V(W_2_29_2) = 1 V(W_2_29_2_bar) = 0
.IC V(W_2_29_3) = 0 V(W_2_29_3_bar) = 1
.IC V(W_2_29_4) = 0 V(W_2_29_4_bar) = 1
.IC V(W_2_30_1) = 1 V(W_2_30_1_bar) = 0
.IC V(W_2_30_2) = 0 V(W_2_30_2_bar) = 1
.IC V(W_2_30_3) = 1 V(W_2_30_3_bar) = 0
.IC V(W_2_30_4) = 0 V(W_2_30_4_bar) = 1
.IC V(W_2_31_1) = 1 V(W_2_31_1_bar) = 0
.IC V(W_2_31_2) = 0 V(W_2_31_2_bar) = 1
.IC V(W_2_31_3) = 1 V(W_2_31_3_bar) = 0
.IC V(W_2_31_4) = 0 V(W_2_31_4_bar) = 1
.IC V(W_2_32_1) = 0 V(W_2_32_1_bar) = 1
.IC V(W_2_32_2) = 1 V(W_2_32_2_bar) = 0
.IC V(W_2_32_3) = 0 V(W_2_32_3_bar) = 1
.IC V(W_2_32_4) = 1 V(W_2_32_4_bar) = 0
.IC V(W_3_1_1) = 1 V(W_3_1_1_bar) = 0
.IC V(W_3_1_2) = 0 V(W_3_1_2_bar) = 1
.IC V(W_3_1_3) = 0 V(W_3_1_3_bar) = 1
.IC V(W_3_1_4) = 1 V(W_3_1_4_bar) = 0
.IC V(W_3_2_1) = 0 V(W_3_2_1_bar) = 1
.IC V(W_3_2_2) = 1 V(W_3_2_2_bar) = 0
.IC V(W_3_2_3) = 1 V(W_3_2_3_bar) = 0
.IC V(W_3_2_4) = 0 V(W_3_2_4_bar) = 1
.IC V(W_3_3_1) = 0 V(W_3_3_1_bar) = 1
.IC V(W_3_3_2) = 1 V(W_3_3_2_bar) = 0
.IC V(W_3_3_3) = 0 V(W_3_3_3_bar) = 1
.IC V(W_3_3_4) = 0 V(W_3_3_4_bar) = 1
.IC V(W_3_4_1) = 1 V(W_3_4_1_bar) = 0
.IC V(W_3_4_2) = 0 V(W_3_4_2_bar) = 1
.IC V(W_3_4_3) = 1 V(W_3_4_3_bar) = 0
.IC V(W_3_4_4) = 0 V(W_3_4_4_bar) = 1
.IC V(W_3_5_1) = 1 V(W_3_5_1_bar) = 0
.IC V(W_3_5_2) = 0 V(W_3_5_2_bar) = 1
.IC V(W_3_5_3) = 0 V(W_3_5_3_bar) = 1
.IC V(W_3_5_4) = 1 V(W_3_5_4_bar) = 0
.IC V(W_3_6_1) = 1 V(W_3_6_1_bar) = 0
.IC V(W_3_6_2) = 0 V(W_3_6_2_bar) = 1
.IC V(W_3_6_3) = 1 V(W_3_6_3_bar) = 0
.IC V(W_3_6_4) = 0 V(W_3_6_4_bar) = 1
.IC V(W_3_7_1) = 0 V(W_3_7_1_bar) = 1
.IC V(W_3_7_2) = 0 V(W_3_7_2_bar) = 1
.IC V(W_3_7_3) = 0 V(W_3_7_3_bar) = 1
.IC V(W_3_7_4) = 1 V(W_3_7_4_bar) = 0
.IC V(W_3_8_1) = 0 V(W_3_8_1_bar) = 1
.IC V(W_3_8_2) = 0 V(W_3_8_2_bar) = 1
.IC V(W_3_8_3) = 0 V(W_3_8_3_bar) = 1
.IC V(W_3_8_4) = 0 V(W_3_8_4_bar) = 1
.IC V(W_3_9_1) = 1 V(W_3_9_1_bar) = 0
.IC V(W_3_9_2) = 1 V(W_3_9_2_bar) = 0
.IC V(W_3_9_3) = 1 V(W_3_9_3_bar) = 0
.IC V(W_3_9_4) = 1 V(W_3_9_4_bar) = 0
.IC V(W_3_10_1) = 1 V(W_3_10_1_bar) = 0
.IC V(W_3_10_2) = 0 V(W_3_10_2_bar) = 1
.IC V(W_3_10_3) = 1 V(W_3_10_3_bar) = 0
.IC V(W_3_10_4) = 1 V(W_3_10_4_bar) = 0
.IC V(W_3_11_1) = 0 V(W_3_11_1_bar) = 1
.IC V(W_3_11_2) = 0 V(W_3_11_2_bar) = 1
.IC V(W_3_11_3) = 1 V(W_3_11_3_bar) = 0
.IC V(W_3_11_4) = 1 V(W_3_11_4_bar) = 0
.IC V(W_3_12_1) = 1 V(W_3_12_1_bar) = 0
.IC V(W_3_12_2) = 1 V(W_3_12_2_bar) = 0
.IC V(W_3_12_3) = 0 V(W_3_12_3_bar) = 1
.IC V(W_3_12_4) = 0 V(W_3_12_4_bar) = 1
.IC V(W_3_13_1) = 1 V(W_3_13_1_bar) = 0
.IC V(W_3_13_2) = 1 V(W_3_13_2_bar) = 0
.IC V(W_3_13_3) = 1 V(W_3_13_3_bar) = 0
.IC V(W_3_13_4) = 0 V(W_3_13_4_bar) = 1
.IC V(W_3_14_1) = 0 V(W_3_14_1_bar) = 1
.IC V(W_3_14_2) = 0 V(W_3_14_2_bar) = 1
.IC V(W_3_14_3) = 0 V(W_3_14_3_bar) = 1
.IC V(W_3_14_4) = 0 V(W_3_14_4_bar) = 1
.IC V(W_3_15_1) = 0 V(W_3_15_1_bar) = 1
.IC V(W_3_15_2) = 1 V(W_3_15_2_bar) = 0
.IC V(W_3_15_3) = 1 V(W_3_15_3_bar) = 0
.IC V(W_3_15_4) = 0 V(W_3_15_4_bar) = 1
.IC V(W_3_16_1) = 0 V(W_3_16_1_bar) = 1
.IC V(W_3_16_2) = 0 V(W_3_16_2_bar) = 1
.IC V(W_3_16_3) = 0 V(W_3_16_3_bar) = 1
.IC V(W_3_16_4) = 0 V(W_3_16_4_bar) = 1
.IC V(W_3_17_1) = 1 V(W_3_17_1_bar) = 0
.IC V(W_3_17_2) = 1 V(W_3_17_2_bar) = 0
.IC V(W_3_17_3) = 1 V(W_3_17_3_bar) = 0
.IC V(W_3_17_4) = 1 V(W_3_17_4_bar) = 0
.IC V(W_3_18_1) = 1 V(W_3_18_1_bar) = 0
.IC V(W_3_18_2) = 0 V(W_3_18_2_bar) = 1
.IC V(W_3_18_3) = 0 V(W_3_18_3_bar) = 1
.IC V(W_3_18_4) = 1 V(W_3_18_4_bar) = 0
.IC V(W_3_19_1) = 1 V(W_3_19_1_bar) = 0
.IC V(W_3_19_2) = 0 V(W_3_19_2_bar) = 1
.IC V(W_3_19_3) = 0 V(W_3_19_3_bar) = 1
.IC V(W_3_19_4) = 0 V(W_3_19_4_bar) = 1
.IC V(W_3_20_1) = 1 V(W_3_20_1_bar) = 0
.IC V(W_3_20_2) = 1 V(W_3_20_2_bar) = 0
.IC V(W_3_20_3) = 0 V(W_3_20_3_bar) = 1
.IC V(W_3_20_4) = 1 V(W_3_20_4_bar) = 0
.IC V(W_3_21_1) = 1 V(W_3_21_1_bar) = 0
.IC V(W_3_21_2) = 1 V(W_3_21_2_bar) = 0
.IC V(W_3_21_3) = 1 V(W_3_21_3_bar) = 0
.IC V(W_3_21_4) = 0 V(W_3_21_4_bar) = 1
.IC V(W_3_22_1) = 0 V(W_3_22_1_bar) = 1
.IC V(W_3_22_2) = 1 V(W_3_22_2_bar) = 0
.IC V(W_3_22_3) = 0 V(W_3_22_3_bar) = 1
.IC V(W_3_22_4) = 1 V(W_3_22_4_bar) = 0
.IC V(W_3_23_1) = 0 V(W_3_23_1_bar) = 1
.IC V(W_3_23_2) = 0 V(W_3_23_2_bar) = 1
.IC V(W_3_23_3) = 0 V(W_3_23_3_bar) = 1
.IC V(W_3_23_4) = 1 V(W_3_23_4_bar) = 0
.IC V(W_3_24_1) = 1 V(W_3_24_1_bar) = 0
.IC V(W_3_24_2) = 1 V(W_3_24_2_bar) = 0
.IC V(W_3_24_3) = 1 V(W_3_24_3_bar) = 0
.IC V(W_3_24_4) = 0 V(W_3_24_4_bar) = 1
.IC V(W_3_25_1) = 1 V(W_3_25_1_bar) = 0
.IC V(W_3_25_2) = 1 V(W_3_25_2_bar) = 0
.IC V(W_3_25_3) = 1 V(W_3_25_3_bar) = 0
.IC V(W_3_25_4) = 0 V(W_3_25_4_bar) = 1
.IC V(W_3_26_1) = 1 V(W_3_26_1_bar) = 0
.IC V(W_3_26_2) = 1 V(W_3_26_2_bar) = 0
.IC V(W_3_26_3) = 1 V(W_3_26_3_bar) = 0
.IC V(W_3_26_4) = 0 V(W_3_26_4_bar) = 1
.IC V(W_3_27_1) = 1 V(W_3_27_1_bar) = 0
.IC V(W_3_27_2) = 1 V(W_3_27_2_bar) = 0
.IC V(W_3_27_3) = 1 V(W_3_27_3_bar) = 0
.IC V(W_3_27_4) = 0 V(W_3_27_4_bar) = 1
.IC V(W_3_28_1) = 1 V(W_3_28_1_bar) = 0
.IC V(W_3_28_2) = 0 V(W_3_28_2_bar) = 1
.IC V(W_3_28_3) = 0 V(W_3_28_3_bar) = 1
.IC V(W_3_28_4) = 0 V(W_3_28_4_bar) = 1
.IC V(W_3_29_1) = 0 V(W_3_29_1_bar) = 1
.IC V(W_3_29_2) = 0 V(W_3_29_2_bar) = 1
.IC V(W_3_29_3) = 0 V(W_3_29_3_bar) = 1
.IC V(W_3_29_4) = 0 V(W_3_29_4_bar) = 1
.IC V(W_3_30_1) = 0 V(W_3_30_1_bar) = 1
.IC V(W_3_30_2) = 0 V(W_3_30_2_bar) = 1
.IC V(W_3_30_3) = 1 V(W_3_30_3_bar) = 0
.IC V(W_3_30_4) = 0 V(W_3_30_4_bar) = 1
.IC V(W_3_31_1) = 1 V(W_3_31_1_bar) = 0
.IC V(W_3_31_2) = 0 V(W_3_31_2_bar) = 1
.IC V(W_3_31_3) = 0 V(W_3_31_3_bar) = 1
.IC V(W_3_31_4) = 1 V(W_3_31_4_bar) = 0
.IC V(W_3_32_1) = 0 V(W_3_32_1_bar) = 1
.IC V(W_3_32_2) = 0 V(W_3_32_2_bar) = 1
.IC V(W_3_32_3) = 1 V(W_3_32_3_bar) = 0
.IC V(W_3_32_4) = 1 V(W_3_32_4_bar) = 0
.IC V(W_4_1_1) = 0 V(W_4_1_1_bar) = 1
.IC V(W_4_1_2) = 1 V(W_4_1_2_bar) = 0
.IC V(W_4_1_3) = 0 V(W_4_1_3_bar) = 1
.IC V(W_4_1_4) = 1 V(W_4_1_4_bar) = 0
.IC V(W_4_2_1) = 1 V(W_4_2_1_bar) = 0
.IC V(W_4_2_2) = 1 V(W_4_2_2_bar) = 0
.IC V(W_4_2_3) = 0 V(W_4_2_3_bar) = 1
.IC V(W_4_2_4) = 1 V(W_4_2_4_bar) = 0
.IC V(W_4_3_1) = 0 V(W_4_3_1_bar) = 1
.IC V(W_4_3_2) = 0 V(W_4_3_2_bar) = 1
.IC V(W_4_3_3) = 1 V(W_4_3_3_bar) = 0
.IC V(W_4_3_4) = 0 V(W_4_3_4_bar) = 1
.IC V(W_4_4_1) = 0 V(W_4_4_1_bar) = 1
.IC V(W_4_4_2) = 0 V(W_4_4_2_bar) = 1
.IC V(W_4_4_3) = 1 V(W_4_4_3_bar) = 0
.IC V(W_4_4_4) = 1 V(W_4_4_4_bar) = 0
.IC V(W_4_5_1) = 1 V(W_4_5_1_bar) = 0
.IC V(W_4_5_2) = 0 V(W_4_5_2_bar) = 1
.IC V(W_4_5_3) = 1 V(W_4_5_3_bar) = 0
.IC V(W_4_5_4) = 0 V(W_4_5_4_bar) = 1
.IC V(W_4_6_1) = 0 V(W_4_6_1_bar) = 1
.IC V(W_4_6_2) = 0 V(W_4_6_2_bar) = 1
.IC V(W_4_6_3) = 1 V(W_4_6_3_bar) = 0
.IC V(W_4_6_4) = 0 V(W_4_6_4_bar) = 1
.IC V(W_4_7_1) = 1 V(W_4_7_1_bar) = 0
.IC V(W_4_7_2) = 0 V(W_4_7_2_bar) = 1
.IC V(W_4_7_3) = 0 V(W_4_7_3_bar) = 1
.IC V(W_4_7_4) = 0 V(W_4_7_4_bar) = 1
.IC V(W_4_8_1) = 0 V(W_4_8_1_bar) = 1
.IC V(W_4_8_2) = 0 V(W_4_8_2_bar) = 1
.IC V(W_4_8_3) = 0 V(W_4_8_3_bar) = 1
.IC V(W_4_8_4) = 0 V(W_4_8_4_bar) = 1
.IC V(W_4_9_1) = 1 V(W_4_9_1_bar) = 0
.IC V(W_4_9_2) = 1 V(W_4_9_2_bar) = 0
.IC V(W_4_9_3) = 1 V(W_4_9_3_bar) = 0
.IC V(W_4_9_4) = 1 V(W_4_9_4_bar) = 0
.IC V(W_4_10_1) = 0 V(W_4_10_1_bar) = 1
.IC V(W_4_10_2) = 0 V(W_4_10_2_bar) = 1
.IC V(W_4_10_3) = 1 V(W_4_10_3_bar) = 0
.IC V(W_4_10_4) = 0 V(W_4_10_4_bar) = 1
.IC V(W_4_11_1) = 1 V(W_4_11_1_bar) = 0
.IC V(W_4_11_2) = 0 V(W_4_11_2_bar) = 1
.IC V(W_4_11_3) = 1 V(W_4_11_3_bar) = 0
.IC V(W_4_11_4) = 1 V(W_4_11_4_bar) = 0
.IC V(W_4_12_1) = 0 V(W_4_12_1_bar) = 1
.IC V(W_4_12_2) = 0 V(W_4_12_2_bar) = 1
.IC V(W_4_12_3) = 1 V(W_4_12_3_bar) = 0
.IC V(W_4_12_4) = 1 V(W_4_12_4_bar) = 0
.IC V(W_4_13_1) = 1 V(W_4_13_1_bar) = 0
.IC V(W_4_13_2) = 0 V(W_4_13_2_bar) = 1
.IC V(W_4_13_3) = 0 V(W_4_13_3_bar) = 1
.IC V(W_4_13_4) = 1 V(W_4_13_4_bar) = 0
.IC V(W_4_14_1) = 0 V(W_4_14_1_bar) = 1
.IC V(W_4_14_2) = 1 V(W_4_14_2_bar) = 0
.IC V(W_4_14_3) = 0 V(W_4_14_3_bar) = 1
.IC V(W_4_14_4) = 1 V(W_4_14_4_bar) = 0
.IC V(W_4_15_1) = 1 V(W_4_15_1_bar) = 0
.IC V(W_4_15_2) = 0 V(W_4_15_2_bar) = 1
.IC V(W_4_15_3) = 0 V(W_4_15_3_bar) = 1
.IC V(W_4_15_4) = 1 V(W_4_15_4_bar) = 0
.IC V(W_4_16_1) = 1 V(W_4_16_1_bar) = 0
.IC V(W_4_16_2) = 0 V(W_4_16_2_bar) = 1
.IC V(W_4_16_3) = 0 V(W_4_16_3_bar) = 1
.IC V(W_4_16_4) = 1 V(W_4_16_4_bar) = 0
.IC V(W_4_17_1) = 0 V(W_4_17_1_bar) = 1
.IC V(W_4_17_2) = 1 V(W_4_17_2_bar) = 0
.IC V(W_4_17_3) = 1 V(W_4_17_3_bar) = 0
.IC V(W_4_17_4) = 1 V(W_4_17_4_bar) = 0
.IC V(W_4_18_1) = 0 V(W_4_18_1_bar) = 1
.IC V(W_4_18_2) = 0 V(W_4_18_2_bar) = 1
.IC V(W_4_18_3) = 0 V(W_4_18_3_bar) = 1
.IC V(W_4_18_4) = 1 V(W_4_18_4_bar) = 0
.IC V(W_4_19_1) = 0 V(W_4_19_1_bar) = 1
.IC V(W_4_19_2) = 0 V(W_4_19_2_bar) = 1
.IC V(W_4_19_3) = 1 V(W_4_19_3_bar) = 0
.IC V(W_4_19_4) = 0 V(W_4_19_4_bar) = 1
.IC V(W_4_20_1) = 0 V(W_4_20_1_bar) = 1
.IC V(W_4_20_2) = 0 V(W_4_20_2_bar) = 1
.IC V(W_4_20_3) = 0 V(W_4_20_3_bar) = 1
.IC V(W_4_20_4) = 0 V(W_4_20_4_bar) = 1
.IC V(W_4_21_1) = 0 V(W_4_21_1_bar) = 1
.IC V(W_4_21_2) = 0 V(W_4_21_2_bar) = 1
.IC V(W_4_21_3) = 0 V(W_4_21_3_bar) = 1
.IC V(W_4_21_4) = 0 V(W_4_21_4_bar) = 1
.IC V(W_4_22_1) = 0 V(W_4_22_1_bar) = 1
.IC V(W_4_22_2) = 1 V(W_4_22_2_bar) = 0
.IC V(W_4_22_3) = 1 V(W_4_22_3_bar) = 0
.IC V(W_4_22_4) = 0 V(W_4_22_4_bar) = 1
.IC V(W_4_23_1) = 1 V(W_4_23_1_bar) = 0
.IC V(W_4_23_2) = 0 V(W_4_23_2_bar) = 1
.IC V(W_4_23_3) = 0 V(W_4_23_3_bar) = 1
.IC V(W_4_23_4) = 0 V(W_4_23_4_bar) = 1
.IC V(W_4_24_1) = 0 V(W_4_24_1_bar) = 1
.IC V(W_4_24_2) = 1 V(W_4_24_2_bar) = 0
.IC V(W_4_24_3) = 0 V(W_4_24_3_bar) = 1
.IC V(W_4_24_4) = 0 V(W_4_24_4_bar) = 1
.IC V(W_4_25_1) = 1 V(W_4_25_1_bar) = 0
.IC V(W_4_25_2) = 0 V(W_4_25_2_bar) = 1
.IC V(W_4_25_3) = 0 V(W_4_25_3_bar) = 1
.IC V(W_4_25_4) = 0 V(W_4_25_4_bar) = 1
.IC V(W_4_26_1) = 1 V(W_4_26_1_bar) = 0
.IC V(W_4_26_2) = 0 V(W_4_26_2_bar) = 1
.IC V(W_4_26_3) = 1 V(W_4_26_3_bar) = 0
.IC V(W_4_26_4) = 1 V(W_4_26_4_bar) = 0
.IC V(W_4_27_1) = 0 V(W_4_27_1_bar) = 1
.IC V(W_4_27_2) = 1 V(W_4_27_2_bar) = 0
.IC V(W_4_27_3) = 1 V(W_4_27_3_bar) = 0
.IC V(W_4_27_4) = 0 V(W_4_27_4_bar) = 1
.IC V(W_4_28_1) = 1 V(W_4_28_1_bar) = 0
.IC V(W_4_28_2) = 1 V(W_4_28_2_bar) = 0
.IC V(W_4_28_3) = 0 V(W_4_28_3_bar) = 1
.IC V(W_4_28_4) = 1 V(W_4_28_4_bar) = 0
.IC V(W_4_29_1) = 0 V(W_4_29_1_bar) = 1
.IC V(W_4_29_2) = 0 V(W_4_29_2_bar) = 1
.IC V(W_4_29_3) = 1 V(W_4_29_3_bar) = 0
.IC V(W_4_29_4) = 1 V(W_4_29_4_bar) = 0
.IC V(W_4_30_1) = 1 V(W_4_30_1_bar) = 0
.IC V(W_4_30_2) = 0 V(W_4_30_2_bar) = 1
.IC V(W_4_30_3) = 1 V(W_4_30_3_bar) = 0
.IC V(W_4_30_4) = 0 V(W_4_30_4_bar) = 1
.IC V(W_4_31_1) = 1 V(W_4_31_1_bar) = 0
.IC V(W_4_31_2) = 1 V(W_4_31_2_bar) = 0
.IC V(W_4_31_3) = 0 V(W_4_31_3_bar) = 1
.IC V(W_4_31_4) = 1 V(W_4_31_4_bar) = 0
.IC V(W_4_32_1) = 1 V(W_4_32_1_bar) = 0
.IC V(W_4_32_2) = 1 V(W_4_32_2_bar) = 0
.IC V(W_4_32_3) = 0 V(W_4_32_3_bar) = 1
.IC V(W_4_32_4) = 1 V(W_4_32_4_bar) = 0

.end
