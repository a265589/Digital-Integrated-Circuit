.SUBCKT Adder_tree VSS VDD  in[127] in[126] in[125] in[124] in[123] in[122] in[121] in[120] in[119] in[118] in[117] in[116] in[115] in[114] in[113] in[112] in[111] in[110] in[109] in[108] in[107] in[106] in[105] in[104] in[103] in[102] in[101] in[100] in[99] in[98] in[97] in[96] in[95] in[94] in[93] in[92] in[91] in[90] in[89] in[88] in[87] in[86] in[85] in[84] in[83] in[82] in[81] in[80] in[79] in[78] in[77] in[76] in[75] in[74] in[73] in[72] in[71] in[70] in[69] in[68] in[67] in[66] in[65] in[64] in[63] in[62] in[61] in[60] in[59] in[58] in[57] in[56] in[55] in[54] in[53] in[52] in[51] in[50] in[49] in[48] in[47] in[46] in[45] in[44] in[43] in[42] in[41] in[40] in[39] in[38] in[37] in[36] in[35] in[34] in[33] in[32] in[31] in[30] in[29] in[28] in[27] in[26] in[25] in[24] in[23] in[22] in[21] in[20] in[19] in[18] in[17] in[16] in[15] in[14] in[13] in[12] in[11] in[10] in[9] in[8] in[7] in[6] in[5] in[4] in[3] in[2] in[1] in[0] out[12] out[11] out[10] out[9] out[8] out[7] out[6] out[5] out[4] out[3] out[2] out[1] out[0]
XDP_OP_94J1_122_9915_U198 VSS VDD  in[4] in[28] in[36] DP_OP_94J1_122_9915_n299 DP_OP_94J1_122_9915_n300 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U197 VSS VDD  in[44] in[52] in[60] DP_OP_94J1_122_9915_n297 DP_OP_94J1_122_9915_n298 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U195 VSS VDD  in[92] in[100] in[108] DP_OP_94J1_122_9915_n293 DP_OP_94J1_122_9915_n294 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U194 VSS VDD  in[116] in[124] in[120] DP_OP_94J1_122_9915_n291 DP_OP_94J1_122_9915_n292 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U193 VSS VDD  in[112] in[104] in[96] DP_OP_94J1_122_9915_n289 DP_OP_94J1_122_9915_n290 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U192 VSS VDD  in[88] in[80] in[72] DP_OP_94J1_122_9915_n287 DP_OP_94J1_122_9915_n288 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U191 VSS VDD  in[64] in[56] in[48] DP_OP_94J1_122_9915_n285 DP_OP_94J1_122_9915_n286 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U186 VSS VDD  DP_OP_94J1_122_9915_n288 DP_OP_94J1_122_9915_n282 DP_OP_94J1_122_9915_n290 DP_OP_94J1_122_9915_n276 DP_OP_94J1_122_9915_n277 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U185 VSS VDD  DP_OP_94J1_122_9915_n292 DP_OP_94J1_122_9915_n294 DP_OP_94J1_122_9915_n296 DP_OP_94J1_122_9915_n274 DP_OP_94J1_122_9915_n275 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U183 VSS VDD  DP_OP_94J1_122_9915_n298 DP_OP_94J1_122_9915_n300 n136 DP_OP_94J1_122_9915_n272 DP_OP_94J1_122_9915_n273 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U180 VSS VDD  in[21] in[29] in[37] DP_OP_94J1_122_9915_n267 DP_OP_94J1_122_9915_n268 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U178 VSS VDD  in[69] in[77] in[85] DP_OP_94J1_122_9915_n263 DP_OP_94J1_122_9915_n264 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U177 VSS VDD  in[93] in[101] in[109] DP_OP_94J1_122_9915_n261 DP_OP_94J1_122_9915_n262 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U174 VSS VDD  in[9] in[65] in[17] DP_OP_94J1_122_9915_n255 DP_OP_94J1_122_9915_n256 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U167 VSS VDD  DP_OP_94J1_122_9915_n243 DP_OP_94J1_122_9915_n295 DP_OP_94J1_122_9915_n283 DP_OP_94J1_122_9915_n244 DP_OP_94J1_122_9915_n245 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U163 VSS VDD  DP_OP_94J1_122_9915_n258 DP_OP_94J1_122_9915_n252 DP_OP_94J1_122_9915_n256 DP_OP_94J1_122_9915_n235 DP_OP_94J1_122_9915_n236 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U162 VSS VDD  DP_OP_94J1_122_9915_n266 DP_OP_94J1_122_9915_n254 DP_OP_94J1_122_9915_n264 DP_OP_94J1_122_9915_n233 DP_OP_94J1_122_9915_n234 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U150 VSS VDD  in[22] in[30] in[38] DP_OP_94J1_122_9915_n215 DP_OP_94J1_122_9915_n216 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U145 VSS VDD  in[94] in[122] in[102] DP_OP_94J1_122_9915_n205 DP_OP_94J1_122_9915_n206 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U143 VSS VDD  in[126] in[50] in[114] DP_OP_94J1_122_9915_n201 DP_OP_94J1_122_9915_n202 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U139 VSS VDD  DP_OP_94J1_122_9915_n265 DP_OP_94J1_122_9915_n194 DP_OP_94J1_122_9915_n267 DP_OP_94J1_122_9915_n195 DP_OP_94J1_122_9915_n196 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U137 VSS VDD  DP_OP_94J1_122_9915_n263 DP_OP_94J1_122_9915_n249 DP_OP_94J1_122_9915_n191 DP_OP_94J1_122_9915_n192 DP_OP_94J1_122_9915_n193 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U136 VSS VDD  DP_OP_94J1_122_9915_n261 DP_OP_94J1_122_9915_n257 DP_OP_94J1_122_9915_n251 DP_OP_94J1_122_9915_n189 DP_OP_94J1_122_9915_n190 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U135 VSS VDD  DP_OP_94J1_122_9915_n259 DP_OP_94J1_122_9915_n253 DP_OP_94J1_122_9915_n255 DP_OP_94J1_122_9915_n187 DP_OP_94J1_122_9915_n188 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U133 VSS VDD  DP_OP_94J1_122_9915_n247 DP_OP_94J1_122_9915_n241 n86 DP_OP_94J1_122_9915_n185 DP_OP_94J1_122_9915_n186 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U130 VSS VDD  DP_OP_94J1_122_9915_n214 DP_OP_94J1_122_9915_n204 DP_OP_94J1_122_9915_n216 DP_OP_94J1_122_9915_n179 DP_OP_94J1_122_9915_n180 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U126 VSS VDD  DP_OP_94J1_122_9915_n190 DP_OP_94J1_122_9915_n188 DP_OP_94J1_122_9915_n193 DP_OP_94J1_122_9915_n172 DP_OP_94J1_122_9915_n173 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U125 VSS VDD  DP_OP_94J1_122_9915_n233 DP_OP_94J1_122_9915_n235 n21 DP_OP_94J1_122_9915_n170 DP_OP_94J1_122_9915_n171 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U121 VSS VDD  DP_OP_94J1_122_9915_n180 DP_OP_94J1_122_9915_n178 n77 DP_OP_94J1_122_9915_n165 DP_OP_94J1_122_9915_n166 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U112 VSS VDD  in[63] in[3] in[71] DP_OP_94J1_122_9915_n149 DP_OP_94J1_122_9915_n150 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U111 VSS VDD  in[79] in[99] in[11] DP_OP_94J1_122_9915_n147 DP_OP_94J1_122_9915_n148 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U110 VSS VDD  in[19] in[107] in[87] DP_OP_94J1_122_9915_n145 DP_OP_94J1_122_9915_n146 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U108 VSS VDD  in[111] in[35] in[119] DP_OP_94J1_122_9915_n141 DP_OP_94J1_122_9915_n142 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U107 VSS VDD  in[127] in[43] in[123] DP_OP_94J1_122_9915_n139 DP_OP_94J1_122_9915_n140 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U106 VSS VDD  in[91] in[51] in[83] DP_OP_94J1_122_9915_n137 DP_OP_94J1_122_9915_n138 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U105 VSS VDD  in[75] in[59] in[67] DP_OP_94J1_122_9915_n135 DP_OP_94J1_122_9915_n136 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U100 VSS VDD  DP_OP_94J1_122_9915_n209 DP_OP_94J1_122_9915_n199 DP_OP_94J1_122_9915_n205 DP_OP_94J1_122_9915_n127 DP_OP_94J1_122_9915_n128 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U99 VSS VDD  DP_OP_94J1_122_9915_n207 DP_OP_94J1_122_9915_n203 DP_OP_94J1_122_9915_n201 DP_OP_94J1_122_9915_n125 DP_OP_94J1_122_9915_n126 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U97 VSS VDD  DP_OP_94J1_122_9915_n189 DP_OP_94J1_122_9915_n195 n14 DP_OP_94J1_122_9915_n123 DP_OP_94J1_122_9915_n124 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U91 VSS VDD  DP_OP_94J1_122_9915_n134 DP_OP_94J1_122_9915_n192 n129 DP_OP_94J1_122_9915_n113 DP_OP_94J1_122_9915_n114 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U89 VSS VDD  DP_OP_94J1_122_9915_n182 DP_OP_94J1_122_9915_n179 n24 DP_OP_94J1_122_9915_n110 DP_OP_94J1_122_9915_n111 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U69 VSS VDD  DP_OP_94J1_122_9915_n137 DP_OP_94J1_122_9915_n151 DP_OP_94J1_122_9915_n149 DP_OP_94J1_122_9915_n80 DP_OP_94J1_122_9915_n81 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U68 VSS VDD  DP_OP_94J1_122_9915_n147 DP_OP_94J1_122_9915_n143 DP_OP_94J1_122_9915_n135 DP_OP_94J1_122_9915_n78 DP_OP_94J1_122_9915_n79 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U67 VSS VDD  DP_OP_94J1_122_9915_n139 DP_OP_94J1_122_9915_n141 DP_OP_94J1_122_9915_n145 DP_OP_94J1_122_9915_n76 DP_OP_94J1_122_9915_n77 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U66 VSS VDD  DP_OP_94J1_122_9915_n130 DP_OP_94J1_122_9915_n133 DP_OP_94J1_122_9915_n125 DP_OP_94J1_122_9915_n74 DP_OP_94J1_122_9915_n75 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U65 VSS VDD  DP_OP_94J1_122_9915_n115 DP_OP_94J1_122_9915_n84 DP_OP_94J1_122_9915_n127 DP_OP_94J1_122_9915_n72 DP_OP_94J1_122_9915_n73 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U62 VSS VDD  DP_OP_94J1_122_9915_n81 DP_OP_94J1_122_9915_n79 DP_OP_94J1_122_9915_n117 DP_OP_94J1_122_9915_n67 DP_OP_94J1_122_9915_n68 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U61 VSS VDD  DP_OP_94J1_122_9915_n75 DP_OP_94J1_122_9915_n113 DP_OP_94J1_122_9915_n107 DP_OP_94J1_122_9915_n65 DP_OP_94J1_122_9915_n66 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U53 VSS VDD  DP_OP_94J1_122_9915_n76 DP_OP_94J1_122_9915_n83 DP_OP_94J1_122_9915_n80 DP_OP_94J1_122_9915_n51 DP_OP_94J1_122_9915_n52 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U51 VSS VDD  DP_OP_94J1_122_9915_n72 DP_OP_94J1_122_9915_n74 n90 DP_OP_94J1_122_9915_n49 DP_OP_94J1_122_9915_n50 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U49 VSS VDD  DP_OP_94J1_122_9915_n63 DP_OP_94J1_122_9915_n65 DP_OP_94J1_122_9915_n50 DP_OP_94J1_122_9915_n44 DP_OP_94J1_122_9915_n45 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U44 VSS VDD  DP_OP_94J1_122_9915_n49 DP_OP_94J1_122_9915_n46 DP_OP_94J1_122_9915_n36 DP_OP_94J1_122_9915_n37 DP_OP_94J1_122_9915_n38 FAx1_ASAP7_75t_R
XDP_OP_94J1_122_9915_U43 VSS VDD  DP_OP_94J1_122_9915_n38 DP_OP_94J1_122_9915_n44 DP_OP_94J1_122_9915_n42 DP_OP_94J1_122_9915_n34 DP_OP_94J1_122_9915_n35 FAx1_ASAP7_75t_R
XU3 VSS VDD  n154 n220 INVx2_ASAP7_75t_R
XU4 VSS VDD  n163 n18 n212 XNOR2xp5_ASAP7_75t_R
XU5 VSS VDD  DP_OP_94J1_122_9915_n90 n6 n132 XNOR2xp5_ASAP7_75t_R
XU6 VSS VDD  n121 n50 n19 XOR2xp5_ASAP7_75t_R
XU7 VSS VDD  n178 n6 BUFx3_ASAP7_75t_R
XU8 VSS VDD  n16 n47 n18 XOR2xp5_ASAP7_75t_R
XU9 VSS VDD  n177 n56 n135 XNOR2xp5_ASAP7_75t_R
XU10 VSS VDD  n130 n71 n121 XNOR2xp5_ASAP7_75t_R
XU11 VSS VDD  n204 n161 DP_OP_94J1_122_9915_n106 XOR2xp5_ASAP7_75t_R
XU12 VSS VDD  DP_OP_94J1_122_9915_n126 DP_OP_94J1_122_9915_n116 n161 XNOR2xp5_ASAP7_75t_R
XU13 VSS VDD  n43 n44 n193 XNOR2xp5_ASAP7_75t_R
XU14 VSS VDD  DP_OP_94J1_122_9915_n131 n158 n54 XNOR2xp5_ASAP7_75t_R
XU15 VSS VDD  DP_OP_94J1_122_9915_n146 n169 n134 XOR2xp5_ASAP7_75t_R
XU16 VSS VDD  DP_OP_94J1_122_9915_n120 DP_OP_94J1_122_9915_n77 n164 XOR2xp5_ASAP7_75t_R
XU17 VSS VDD  DP_OP_94J1_122_9915_n170 n168 n167 XNOR2xp5_ASAP7_75t_R
XU18 VSS VDD  DP_OP_94J1_122_9915_n48 n90 INVx3_ASAP7_75t_R
XU19 VSS VDD  DP_OP_94J1_122_9915_n177 n89 n158 XNOR2xp5_ASAP7_75t_R
XU20 VSS VDD  n26 n180 n93 XOR2xp5_ASAP7_75t_R
XU21 VSS VDD  n40 n148 INVx1_ASAP7_75t_R
XU22 VSS VDD  n33 n173 INVx1_ASAP7_75t_R
XU23 VSS VDD  n13 n12 DP_OP_94J1_122_9915_n121 XOR2x2_ASAP7_75t_R
XU24 VSS VDD  in[23] n205 DP_OP_94J1_122_9915_n154 XNOR2x2_ASAP7_75t_R
XU25 VSS VDD  n153 n184 DP_OP_94J1_122_9915_n240 XNOR2xp5_ASAP7_75t_R
XU26 VSS VDD  in[7] in[15] DP_OP_94J1_122_9915_n129 XNOR2xp5_ASAP7_75t_R
XU27 VSS VDD  in[117] in[1] n181 XNOR2xp5_ASAP7_75t_R
XU28 VSS VDD  in[57] in[49] n183 XNOR2xp5_ASAP7_75t_R
XU29 VSS VDD  in[13] in[5] DP_OP_94J1_122_9915_n194 NAND2xp5_ASAP7_75t_R
XU30 VSS VDD  n5 TIEHIx1_ASAP7_75t_R
XU31 VSS VDD  n5 out[9] INVx1_ASAP7_75t_R
XU32 VSS VDD  n5 out[10] INVx1_ASAP7_75t_R
XU33 VSS VDD  n5 out[11] INVx1_ASAP7_75t_R
XU34 VSS VDD  n5 out[12] INVx1_ASAP7_75t_R
XU35 VSS VDD  n62 n219 out[6] XNOR2xp5_ASAP7_75t_R
XU36 VSS VDD  n56 n126 n123 NAND2xp5_ASAP7_75t_R
XU37 VSS VDD  n36 n149 n165 XNOR2x1_ASAP7_75t_R
XU38 VSS VDD  DP_OP_94J1_122_9915_n185 n24 INVx1_ASAP7_75t_R
XU39 VSS VDD  n121 n50 n22 XNOR2xp5_ASAP7_75t_R
XU40 VSS VDD  n7 DP_OP_94J1_122_9915_n63 n99 XOR2xp5_ASAP7_75t_R
XU41 VSS VDD  DP_OP_94J1_122_9915_n65 n8 n7 XOR2xp5_ASAP7_75t_R
XU42 VSS VDD  DP_OP_94J1_122_9915_n50 n8 INVx1_ASAP7_75t_R
XU43 VSS VDD  DP_OP_94J1_122_9915_n196 n202 DP_OP_94J1_122_9915_n176 XOR2xp5_ASAP7_75t_R
XU44 VSS VDD  in[14] in[6] DP_OP_94J1_122_9915_n191 XNOR2xp5_ASAP7_75t_R
XU45 VSS VDD  n40 n33 n84 NAND2xp5_ASAP7_75t_R
XU46 VSS VDD  n9 n215 out[4] XOR2xp5_ASAP7_75t_R
XU47 VSS VDD  DP_OP_94J1_122_9915_n57 n216 n9 XOR2xp5_ASAP7_75t_R
XU48 VSS VDD  n10 n178 n131 XNOR2xp5_ASAP7_75t_R
XU49 VSS VDD  n35 n177 n178 XNOR2x1_ASAP7_75t_R
XU50 VSS VDD  n48 n49 DP_OP_94J1_122_9915_n284 XNOR2x1_ASAP7_75t_R
XU51 VSS VDD  n98 n25 n110 NAND2xp5_ASAP7_75t_R
XU52 VSS VDD  DP_OP_94J1_122_9915_n272 n25 INVx1_ASAP7_75t_R
XU53 VSS VDD  n115 n114 n10 NAND2xp5_ASAP7_75t_R
XU54 VSS VDD  n15 DP_OP_94J1_122_9915_n172 DP_OP_94J1_122_9915_n114 DP_OP_94J1_122_9915_n99 MAJIxp5_ASAP7_75t_R
XU55 VSS VDD  n11 n15 DP_OP_94J1_122_9915_n100 XNOR2xp5_ASAP7_75t_R
XU56 VSS VDD  DP_OP_94J1_122_9915_n114 DP_OP_94J1_122_9915_n172 n11 XOR2xp5_ASAP7_75t_R
XU57 VSS VDD  n13 DP_OP_94J1_122_9915_n136 DP_OP_94J1_122_9915_n150 DP_OP_94J1_122_9915_n120 MAJIxp5_ASAP7_75t_R
XU58 VSS VDD  DP_OP_94J1_122_9915_n136 DP_OP_94J1_122_9915_n150 n12 XNOR2xp5_ASAP7_75t_R
XU59 VSS VDD  DP_OP_94J1_122_9915_n187 n13 INVx1_ASAP7_75t_R
XU60 VSS VDD  DP_OP_94J1_122_9915_n140 n137 BUFx2_ASAP7_75t_R
XU61 VSS VDD  n137 n14 INVx2_ASAP7_75t_R
XU62 VSS VDD  DP_OP_94J1_122_9915_n121 n15 INVx2_ASAP7_75t_R
XU63 VSS VDD  DP_OP_94J1_122_9915_n245 DP_OP_94J1_122_9915_n240 DP_OP_94J1_122_9915_n242 n16 MAJIxp5_ASAP7_75t_R
XU64 VSS VDD  DP_OP_94J1_122_9915_n243 DP_OP_94J1_122_9915_n283 DP_OP_94J1_122_9915_n295 A0  n17 FAx1_ASAP7_75t_R
XU65 VSS VDD  n38 n45 INVx2_ASAP7_75t_R
XU66 VSS VDD  n42 n45 DP_OP_94J1_122_9915_n97 XNOR2x2_ASAP7_75t_R
XU67 VSS VDD  DP_OP_94J1_122_9915_n97 n64 n127 XNOR2xp5_ASAP7_75t_R
XU68 VSS VDD  n217 n19 n218 XNOR2xp5_ASAP7_75t_R
XU69 VSS VDD  n135 DP_OP_94J1_122_9915_n90 n195 n20 MAJIxp5_ASAP7_75t_R
XU70 VSS VDD  n195 DP_OP_94J1_122_9915_n90 n135 n217 MAJx2_ASAP7_75t_R
XU71 VSS VDD  DP_OP_94J1_122_9915_n262 n144 n145 n21 MAJIxp5_ASAP7_75t_R
XU72 VSS VDD  n16 n47 n23 XNOR2xp5_ASAP7_75t_R
XU73 VSS VDD  in[93] in[101] in[109] A1  n26 FAx1_ASAP7_75t_R
XU74 VSS VDD  in[94] in[122] in[102] n27 MAJIxp5_ASAP7_75t_R
XU75 VSS VDD  DP_OP_94J1_122_9915_n173 n172 n108 NAND2xp5_ASAP7_75t_R
XU76 VSS VDD  DP_OP_94J1_122_9915_n221 n193 n163 XNOR2xp5_ASAP7_75t_R
XU77 VSS VDD  in[44] in[52] in[60] n28 MAJIxp5_ASAP7_75t_R
XU78 VSS VDD  n51 n20 n22 n219 MAJx2_ASAP7_75t_R
XU79 VSS VDD  DP_OP_94J1_122_9915_n111 n38 BUFx4_ASAP7_75t_R
XU80 VSS VDD  DP_OP_94J1_122_9915_n166 n100 BUFx4_ASAP7_75t_R
XU81 VSS VDD  DP_OP_94J1_122_9915_n78 DP_OP_94J1_122_9915_n48 BUFx5_ASAP7_75t_R
XU82 VSS VDD  n138 n77 INVx3_ASAP7_75t_R
XU83 VSS VDD  in[40] n49 INVx8_ASAP7_75t_R
XU84 VSS VDD  n147 n170 INVx3_ASAP7_75t_R
XU85 VSS VDD  DP_OP_94J1_122_9915_n236 n33 BUFx4_ASAP7_75t_R
XU86 VSS VDD  DP_OP_94J1_122_9915_n234 n40 BUFx4_ASAP7_75t_R
XU87 VSS VDD  DP_OP_94J1_122_9915_n124 n147 BUFx4_ASAP7_75t_R
XU88 VSS VDD  DP_OP_94J1_122_9915_n66 n56 BUFx4_ASAP7_75t_R
XU89 VSS VDD  in[20] in[12] n29 AND2x2_ASAP7_75t_R
XU90 VSS VDD  n204 n161 n30 XNOR2xp5_ASAP7_75t_R
XU91 VSS VDD  in[86] n57 n31 XOR2xp5_ASAP7_75t_R
XU92 VSS VDD  DP_OP_94J1_122_9915_n62 DP_OP_94J1_122_9915_n93 DP_OP_94J1_122_9915_n64 n32 MAJx2_ASAP7_75t_R
XU93 VSS VDD  n56 n35 INVx3_ASAP7_75t_R
XU94 VSS VDD  DP_OP_94J1_122_9915_n186 n138 BUFx4_ASAP7_75t_R
XU95 VSS VDD  DP_OP_94J1_122_9915_n180 DP_OP_94J1_122_9915_n178 n77 n36 MAJx2_ASAP7_75t_R
XU96 VSS VDD  in[20] in[12] n34 NAND2xp33_ASAP7_75t_R
XU97 VSS VDD  DP_OP_94J1_122_9915_n69 n78 INVx4_ASAP7_75t_R
XU98 VSS VDD  DP_OP_94J1_122_9915_n123 DP_OP_94J1_122_9915_n69 BUFx5_ASAP7_75t_R
XU99 VSS VDD  DP_OP_94J1_122_9915_n298 DP_OP_94J1_122_9915_n300 n136 n37 MAJIxp5_ASAP7_75t_R
XU100 VSS VDD  DP_OP_94J1_122_9915_n62 DP_OP_94J1_122_9915_n93 DP_OP_94J1_122_9915_n64 n39 MAJIxp5_ASAP7_75t_R
XU101 VSS VDD  DP_OP_94J1_122_9915_n128 n89 INVx1_ASAP7_75t_R
XU102 VSS VDD  n31 DP_OP_94J1_122_9915_n244 DP_OP_94J1_122_9915_n196 n204 MAJx2_ASAP7_75t_R
XU103 VSS VDD  in[32] in[0] n48 XNOR2xp5_ASAP7_75t_R
XU104 VSS VDD  DP_OP_94J1_122_9915_n232 n84 n117 NAND2xp33_ASAP7_75t_R
XU105 VSS VDD  DP_OP_94J1_122_9915_n245 n201 n98 XOR2xp5_ASAP7_75t_R
XU106 VSS VDD  n100 n106 INVx1_ASAP7_75t_R
XU107 VSS VDD  n167 n170 n97 XOR2xp5_ASAP7_75t_R
XU108 VSS VDD  n167 n170 n83 XNOR2xp5_ASAP7_75t_R
XU109 VSS VDD  DP_OP_94J1_122_9915_n226 DP_OP_94J1_122_9915_n176 n44 XNOR2xp5_ASAP7_75t_R
XU110 VSS VDD  n148 n173 n118 NAND2xp33_ASAP7_75t_R
XU111 VSS VDD  DP_OP_94J1_122_9915_n248 n111 DP_OP_94J1_122_9915_n232 XOR2xp5_ASAP7_75t_R
XU112 VSS VDD  n93 n186 n94 XNOR2xp5_ASAP7_75t_R
XU113 VSS VDD  in[7] in[15] n221 NAND2xp5_ASAP7_75t_R
XU114 VSS VDD  in[68] in[84] in[76] DP_OP_94J1_122_9915_n295 MAJIxp5_ASAP7_75t_R
XU115 VSS VDD  in[68] n41 DP_OP_94J1_122_9915_n296 XNOR2xp5_ASAP7_75t_R
XU116 VSS VDD  in[84] in[76] n41 XOR2xp5_ASAP7_75t_R
XU117 VSS VDD  n103 n54 n42 XNOR2xp5_ASAP7_75t_R
XU118 VSS VDD  n65 DP_OP_94J1_122_9915_n231 n87 n103 MAJx2_ASAP7_75t_R
XU119 VSS VDD  DP_OP_94J1_122_9915_n97 n64 n69 XOR2xp5_ASAP7_75t_R
XU120 VSS VDD  DP_OP_94J1_122_9915_n221 n23 n193 n64 MAJx2_ASAP7_75t_R
XU121 VSS VDD  n55 n46 DP_OP_94J1_122_9915_n221 NAND2xp5_ASAP7_75t_R
XU122 VSS VDD  n95 n43 INVx1_ASAP7_75t_R
XU123 VSS VDD  n81 n110 n46 NAND2xp5_ASAP7_75t_R
XU124 VSS VDD  DP_OP_94J1_122_9915_n231 n87 n47 XOR2xp5_ASAP7_75t_R
XU125 VSS VDD  DP_OP_94J1_122_9915_n278 DP_OP_94J1_122_9915_n284 n171 XNOR2xp5_ASAP7_75t_R
XU126 VSS VDD  n32 n52 n50 XNOR2xp5_ASAP7_75t_R
XU127 VSS VDD  n140 DP_OP_94J1_122_9915_n57 n216 n51 MAJIxp5_ASAP7_75t_R
XU128 VSS VDD  n67 DP_OP_94J1_122_9915_n91 n68 n216 MAJx2_ASAP7_75t_R
XU129 VSS VDD  n195 n131 n140 XNOR2xp5_ASAP7_75t_R
XU130 VSS VDD  n219 DP_OP_94J1_122_9915_n39 DP_OP_94J1_122_9915_n35 n53 MAJIxp5_ASAP7_75t_R
XU131 VSS VDD  n99 n52 INVxp67_ASAP7_75t_R
XU132 VSS VDD  n223 n53 out[7] XNOR2xp5_ASAP7_75t_R
XU133 VSS VDD  n220 DP_OP_94J1_122_9915_n37 n53 out[8] MAJIxp5_ASAP7_75t_R
XU134 VSS VDD  n37 n80 n55 NAND2xp33_ASAP7_75t_R
XU135 VSS VDD  n35 n125 n124 NAND2xp33_ASAP7_75t_R
XU136 VSS VDD  in[86] in[34] in[26] DP_OP_94J1_122_9915_n207 MAJIxp5_ASAP7_75t_R
XU137 VSS VDD  in[34] in[26] n57 XOR2xp5_ASAP7_75t_R
XU138 VSS VDD  DP_OP_94J1_122_9915_n144 DP_OP_94J1_122_9915_n154 n58 DP_OP_94J1_122_9915_n115 MAJIxp5_ASAP7_75t_R
XU139 VSS VDD  n59 n58 DP_OP_94J1_122_9915_n116 XNOR2xp5_ASAP7_75t_R
XU140 VSS VDD  in[47] n200 n58 XNOR2xp5_ASAP7_75t_R
XU141 VSS VDD  DP_OP_94J1_122_9915_n144 DP_OP_94J1_122_9915_n154 n59 XOR2xp5_ASAP7_75t_R
XU142 VSS VDD  n60 n109 n108 n114 NAND3xp33_ASAP7_75t_R
XU143 VSS VDD  n60 n113 DP_OP_94J1_122_9915_n90 NAND2xp5_ASAP7_75t_R
XU144 VSS VDD  n107 n83 n60 NAND2xp5_ASAP7_75t_R
XU145 VSS VDD  DP_OP_94J1_122_9915_n206 DP_OP_94J1_122_9915_n200 DP_OP_94J1_122_9915_n212 DP_OP_94J1_122_9915_n177 MAJIxp5_ASAP7_75t_R
XU146 VSS VDD  n61 DP_OP_94J1_122_9915_n206 DP_OP_94J1_122_9915_n178 XOR2xp5_ASAP7_75t_R
XU147 VSS VDD  DP_OP_94J1_122_9915_n200 DP_OP_94J1_122_9915_n212 n61 XNOR2xp5_ASAP7_75t_R
XU148 VSS VDD  DP_OP_94J1_122_9915_n39 DP_OP_94J1_122_9915_n35 n62 XNOR2xp5_ASAP7_75t_R
XU149 VSS VDD  n120 n63 DP_OP_94J1_122_9915_n39 NAND2xp5_ASAP7_75t_R
XU150 VSS VDD  n121 n119 n63 NAND2xp5_ASAP7_75t_R
XU151 VSS VDD  DP_OP_94J1_122_9915_n94 DP_OP_94J1_122_9915_n97 n64 n195 MAJIxp5_ASAP7_75t_R
XU152 VSS VDD  n17 DP_OP_94J1_122_9915_n240 DP_OP_94J1_122_9915_n242 n65 MAJIxp5_ASAP7_75t_R
XU153 VSS VDD  n34 DP_OP_94J1_122_9915_n297 DP_OP_94J1_122_9915_n299 DP_OP_94J1_122_9915_n247 MAJIxp5_ASAP7_75t_R
XU154 VSS VDD  n28 n66 DP_OP_94J1_122_9915_n248 XNOR2xp5_ASAP7_75t_R
XU155 VSS VDD  n29 DP_OP_94J1_122_9915_n299 n66 XNOR2xp5_ASAP7_75t_R
XU156 VSS VDD  n142 DP_OP_94J1_122_9915_n161 n188 n67 MAJIxp5_ASAP7_75t_R
XU157 VSS VDD  n163 n23 n142 XNOR2xp5_ASAP7_75t_R
XU158 VSS VDD  n72 n69 n68 XNOR2xp5_ASAP7_75t_R
XU159 VSS VDD  n30 n165 n72 XOR2xp5_ASAP7_75t_R
XU160 VSS VDD  n100 n70 DP_OP_94J1_122_9915_n161 XOR2x2_ASAP7_75t_R
XU161 VSS VDD  DP_OP_94J1_122_9915_n173 n172 n70 XNOR2xp5_ASAP7_75t_R
XU162 VSS VDD  n126 n124 n71 NAND2xp5_ASAP7_75t_R
XU163 VSS VDD  n142 n188 DP_OP_94J1_122_9915_n161 n73 MAJIxp5_ASAP7_75t_R
XU164 VSS VDD  in[58] in[66] in[90] n74 MAJIxp5_ASAP7_75t_R
XU165 VSS VDD  DP_OP_94J1_122_9915_n99 DP_OP_94J1_122_9915_n96 n177 XOR2x2_ASAP7_75t_R
XU166 VSS VDD  in[25] in[97] n206 XOR2xp5_ASAP7_75t_R
XU167 VSS VDD  in[66] in[90] n207 XOR2xp5_ASAP7_75t_R
XU168 VSS VDD  DP_OP_94J1_122_9915_n274 DP_OP_94J1_122_9915_n276 n186 XNOR2xp5_ASAP7_75t_R
XU169 VSS VDD  DP_OP_94J1_122_9915_n106 n165 DP_OP_94J1_122_9915_n94 XNOR2xp5_ASAP7_75t_R
XU170 VSS VDD  in[73] in[33] n203 XOR2xp5_ASAP7_75t_R
XU171 VSS VDD  in[118] in[42] n190 XOR2xp5_ASAP7_75t_R
XU172 VSS VDD  in[55] in[115] n200 XOR2xp5_ASAP7_75t_R
XU173 VSS VDD  in[81] n181 n146 XNOR2xp5_ASAP7_75t_R
XU174 VSS VDD  DP_OP_94J1_122_9915_n210 DP_OP_94J1_122_9915_n202 n101 XNOR2xp5_ASAP7_75t_R
XU175 VSS VDD  in[61] in[53] n192 XOR2xp5_ASAP7_75t_R
XU176 VSS VDD  in[10] in[106] n191 XOR2xp5_ASAP7_75t_R
XU177 VSS VDD  in[20] in[12] DP_OP_94J1_122_9915_n278 XNOR2xp5_ASAP7_75t_R
XU178 VSS VDD  in[16] in[8] n199 XOR2xp5_ASAP7_75t_R
XU179 VSS VDD  n194 n82 n209 XNOR2xp5_ASAP7_75t_R
XU180 VSS VDD  DP_OP_94J1_122_9915_n45 n39 n119 NAND2xp33_ASAP7_75t_R
XU181 VSS VDD  n128 DP_OP_94J1_122_9915_n91 n214 XOR2xp5_ASAP7_75t_R
XU182 VSS VDD  n78 DP_OP_94J1_122_9915_n77 DP_OP_94J1_122_9915_n120 n76 MAJIxp5_ASAP7_75t_R
XU183 VSS VDD  n78 DP_OP_94J1_122_9915_n77 DP_OP_94J1_122_9915_n120 DP_OP_94J1_122_9915_n70 MAJx2_ASAP7_75t_R
XU184 VSS VDD  n92 n105 n79 NAND2xp5_ASAP7_75t_R
XU185 VSS VDD  n17 n201 n80 XNOR2xp5_ASAP7_75t_R
XU186 VSS VDD  n93 n186 n81 XOR2xp5_ASAP7_75t_R
XU187 VSS VDD  n111 DP_OP_94J1_122_9915_n248 n82 XNOR2xp5_ASAP7_75t_R
XU188 VSS VDD  in[106] in[10] in[2] n85 MAJIxp5_ASAP7_75t_R
XU189 VSS VDD  in[74] n116 n86 XOR2xp5_ASAP7_75t_R
XU190 VSS VDD  n102 n101 n87 XNOR2xp5_ASAP7_75t_R
XU191 VSS VDD  n105 n92 n88 AND2x2_ASAP7_75t_R
XU192 VSS VDD  n39 DP_OP_94J1_122_9915_n45 n120 OR2x2_ASAP7_75t_R
XU193 VSS VDD  in[106] in[10] in[2] n91 MAJx2_ASAP7_75t_R
XU194 VSS VDD  DP_OP_94J1_122_9915_n173 n172 n92 OR2x2_ASAP7_75t_R
XU195 VSS VDD  DP_OP_94J1_122_9915_n99 DP_OP_94J1_122_9915_n96 n125 NAND2xp33_ASAP7_75t_R
XU196 VSS VDD  n100 n92 n109 NAND2xp33_ASAP7_75t_R
XU197 VSS VDD  DP_OP_94J1_122_9915_n233 n21 DP_OP_94J1_122_9915_n235 n75 n95 FAx1_ASAP7_75t_R
XU198 VSS VDD  DP_OP_94J1_122_9915_n209 n74 n27 A2  n96 FAx1_ASAP7_75t_R
XU199 VSS VDD  DP_OP_94J1_122_9915_n202 DP_OP_94J1_122_9915_n210 n102 DP_OP_94J1_122_9915_n182 MAJIxp5_ASAP7_75t_R
XU200 VSS VDD  DP_OP_94J1_122_9915_n293 DP_OP_94J1_122_9915_n289 DP_OP_94J1_122_9915_n291 n102 MAJx2_ASAP7_75t_R
XU201 VSS VDD  n38 n104 n103 DP_OP_94J1_122_9915_n96 MAJIxp5_ASAP7_75t_R
XU202 VSS VDD  DP_OP_94J1_122_9915_n131 n158 n104 XNOR2xp5_ASAP7_75t_R
XU203 VSS VDD  n106 n108 n105 NAND2xp5_ASAP7_75t_R
XU204 VSS VDD  DP_OP_94J1_122_9915_n100 n107 INVx1_ASAP7_75t_R
XU205 VSS VDD  DP_OP_94J1_122_9915_n230 n112 DP_OP_94J1_122_9915_n248 DP_OP_94J1_122_9915_n231 MAJIxp5_ASAP7_75t_R
XU206 VSS VDD  n112 DP_OP_94J1_122_9915_n230 n111 XNOR2xp5_ASAP7_75t_R
XU207 VSS VDD  DP_OP_94J1_122_9915_n286 DP_OP_94J1_122_9915_n284 DP_OP_94J1_122_9915_n278 n112 MAJIxp5_ASAP7_75t_R
XU208 VSS VDD  n115 n88 n113 NAND2xp5_ASAP7_75t_R
XU209 VSS VDD  DP_OP_94J1_122_9915_n100 n97 n115 NAND2xp33_ASAP7_75t_R
XU210 VSS VDD  in[98] in[82] n116 XOR2xp5_ASAP7_75t_R
XU211 VSS VDD  n118 n117 n172 NAND2xp5_ASAP7_75t_R
XU212 VSS VDD  n85 DP_OP_94J1_122_9915_n197 DP_OP_94J1_122_9915_n129 DP_OP_94J1_122_9915_n130 MAJIxp5_ASAP7_75t_R
XU213 VSS VDD  n91 n122 DP_OP_94J1_122_9915_n131 XNOR2xp5_ASAP7_75t_R
XU214 VSS VDD  DP_OP_94J1_122_9915_n129 DP_OP_94J1_122_9915_n197 n122 XNOR2xp5_ASAP7_75t_R
XU215 VSS VDD  in[98] in[82] in[74] DP_OP_94J1_122_9915_n197 MAJIxp5_ASAP7_75t_R
XU216 VSS VDD  n196 n125 n123 n197 NAND3xp33_ASAP7_75t_R
XU217 VSS VDD  DP_OP_94J1_122_9915_n99 DP_OP_94J1_122_9915_n96 n126 OR2x2_ASAP7_75t_R
XU218 VSS VDD  n72 n127 n128 XOR2xp5_ASAP7_75t_R
XU219 VSS VDD  DP_OP_94J1_122_9915_n138 DP_OP_94J1_122_9915_n112 BUFx2_ASAP7_75t_R
XU220 VSS VDD  DP_OP_94J1_122_9915_n112 n129 INVx2_ASAP7_75t_R
XU221 VSS VDD  DP_OP_94J1_122_9915_n47 DP_OP_94J1_122_9915_n61 n130 XOR2xp5_ASAP7_75t_R
XU222 VSS VDD  n198 n197 DP_OP_94J1_122_9915_n42 NAND2xp5_ASAP7_75t_R
XU223 VSS VDD  n195 n132 n215 XNOR2xp5_ASAP7_75t_R
XU224 VSS VDD  n94 n187 n133 XOR2xp5_ASAP7_75t_R
XU225 VSS VDD  DP_OP_94J1_122_9915_n286 n171 n136 XNOR2xp5_ASAP7_75t_R
XU226 VSS VDD  n94 n187 DP_OP_94J1_122_9915_n222 XNOR2xp5_ASAP7_75t_R
XU227 VSS VDD  DP_OP_94J1_122_9915_n146 n169 n168 XNOR2xp5_ASAP7_75t_R
XU228 VSS VDD  in[22] in[30] in[38] n141 MAJIxp5_ASAP7_75t_R
XU229 VSS VDD  n140 DP_OP_94J1_122_9915_n57 n216 n143 MAJIxp5_ASAP7_75t_R
XU230 VSS VDD  DP_OP_94J1_122_9915_n171 DP_OP_94J1_122_9915_n226 DP_OP_94J1_122_9915_n176 n149 MAJx2_ASAP7_75t_R
XU231 VSS VDD  in[41] n183 n144 XOR2xp5_ASAP7_75t_R
XU232 VSS VDD  in[81] n181 n145 XOR2xp5_ASAP7_75t_R
XU233 VSS VDD  DP_OP_94J1_122_9915_n34 n154 BUFx5_ASAP7_75t_R
XU234 VSS VDD  n147 n134 n75 n150 MAJx2_ASAP7_75t_R
XU235 VSS VDD  in[92] in[100] in[108] n153 MAJx2_ASAP7_75t_R
XU236 VSS VDD  in[46] in[62] in[54] n151 MAJx2_ASAP7_75t_R
XU237 VSS VDD  in[88] in[80] in[72] n152 MAJx2_ASAP7_75t_R
XU238 VSS VDD  n33 n40 n194 XOR2x2_ASAP7_75t_R
XU239 VSS VDD  DP_OP_94J1_122_9915_n268 DP_OP_94J1_122_9915_n230 INVx1_ASAP7_75t_R
XU240 VSS VDD  n79 n185 DP_OP_94J1_122_9915_n91 XOR2x2_ASAP7_75t_R
XU241 VSS VDD  DP_OP_94J1_122_9915_n110 DP_OP_94J1_122_9915_n73 n156 DP_OP_94J1_122_9915_n63 MAJIxp5_ASAP7_75t_R
XU242 VSS VDD  n156 n155 DP_OP_94J1_122_9915_n64 XOR2xp5_ASAP7_75t_R
XU243 VSS VDD  DP_OP_94J1_122_9915_n110 DP_OP_94J1_122_9915_n73 n155 XNOR2xp5_ASAP7_75t_R
XU244 VSS VDD  n204 DP_OP_94J1_122_9915_n116 DP_OP_94J1_122_9915_n126 n156 MAJIxp5_ASAP7_75t_R
XU245 VSS VDD  in[13] in[5] DP_OP_94J1_122_9915_n243 XNOR2xp5_ASAP7_75t_R
XU246 VSS VDD  in[46] in[62] in[54] DP_OP_94J1_122_9915_n213 MAJIxp5_ASAP7_75t_R
XU247 VSS VDD  in[46] n157 DP_OP_94J1_122_9915_n214 XNOR2xp5_ASAP7_75t_R
XU248 VSS VDD  in[62] in[54] n157 XOR2xp5_ASAP7_75t_R
XU249 VSS VDD  DP_OP_94J1_122_9915_n131 DP_OP_94J1_122_9915_n177 n96 DP_OP_94J1_122_9915_n107 MAJIxp5_ASAP7_75t_R
XU250 VSS VDD  DP_OP_94J1_122_9915_n287 DP_OP_94J1_122_9915_n281 DP_OP_94J1_122_9915_n285 DP_OP_94J1_122_9915_n241 MAJIxp5_ASAP7_75t_R
XU251 VSS VDD  DP_OP_94J1_122_9915_n242 DP_OP_94J1_122_9915_n240 n201 XNOR2xp5_ASAP7_75t_R
XU252 VSS VDD  n152 n159 DP_OP_94J1_122_9915_n242 XNOR2xp5_ASAP7_75t_R
XU253 VSS VDD  DP_OP_94J1_122_9915_n281 DP_OP_94J1_122_9915_n285 n159 XNOR2xp5_ASAP7_75t_R
XU254 VSS VDD  n76 DP_OP_94J1_122_9915_n52 DP_OP_94J1_122_9915_n67 DP_OP_94J1_122_9915_n46 MAJIxp5_ASAP7_75t_R
XU255 VSS VDD  n160 DP_OP_94J1_122_9915_n70 DP_OP_94J1_122_9915_n47 XNOR2xp5_ASAP7_75t_R
XU256 VSS VDD  DP_OP_94J1_122_9915_n52 DP_OP_94J1_122_9915_n67 n160 XNOR2xp5_ASAP7_75t_R
XU257 VSS VDD  in[40] in[32] in[0] DP_OP_94J1_122_9915_n283 MAJIxp5_ASAP7_75t_R
XU258 VSS VDD  in[95] in[103] in[27] DP_OP_94J1_122_9915_n143 MAJIxp5_ASAP7_75t_R
XU259 VSS VDD  in[95] n162 DP_OP_94J1_122_9915_n144 XNOR2xp5_ASAP7_75t_R
XU260 VSS VDD  in[103] in[27] n162 XOR2xp5_ASAP7_75t_R
XU261 VSS VDD  n164 n78 DP_OP_94J1_122_9915_n71 XNOR2xp5_ASAP7_75t_R
XU262 VSS VDD  DP_OP_94J1_122_9915_n165 DP_OP_94J1_122_9915_n106 n149 DP_OP_94J1_122_9915_n93 MAJIxp5_ASAP7_75t_R
XU263 VSS VDD  DP_OP_94J1_122_9915_n71 n150 DP_OP_94J1_122_9915_n68 DP_OP_94J1_122_9915_n61 MAJIxp5_ASAP7_75t_R
XU264 VSS VDD  DP_OP_94J1_122_9915_n71 n166 DP_OP_94J1_122_9915_n62 XOR2xp5_ASAP7_75t_R
XU265 VSS VDD  DP_OP_94J1_122_9915_n68 n150 n166 XNOR2xp5_ASAP7_75t_R
XU266 VSS VDD  DP_OP_94J1_122_9915_n148 DP_OP_94J1_122_9915_n142 n169 XOR2xp5_ASAP7_75t_R
XU267 VSS VDD  in[70] in[78] in[18] DP_OP_94J1_122_9915_n209 MAJIxp5_ASAP7_75t_R
XU268 VSS VDD  in[70] n174 DP_OP_94J1_122_9915_n210 XNOR2xp5_ASAP7_75t_R
XU269 VSS VDD  in[78] in[18] n174 XOR2xp5_ASAP7_75t_R
XU270 VSS VDD  DP_OP_94J1_122_9915_n213 n176 n141 DP_OP_94J1_122_9915_n133 MAJIxp5_ASAP7_75t_R
XU271 VSS VDD  n151 n175 DP_OP_94J1_122_9915_n134 XNOR2xp5_ASAP7_75t_R
XU272 VSS VDD  n176 DP_OP_94J1_122_9915_n215 n175 XNOR2xp5_ASAP7_75t_R
XU273 VSS VDD  in[6] in[14] n176 NAND2xp5_ASAP7_75t_R
XU274 VSS VDD  in[125] in[121] in[89] DP_OP_94J1_122_9915_n257 MAJIxp5_ASAP7_75t_R
XU275 VSS VDD  in[125] n179 DP_OP_94J1_122_9915_n258 XNOR2xp5_ASAP7_75t_R
XU276 VSS VDD  in[121] in[89] n179 XOR2xp5_ASAP7_75t_R
XU277 VSS VDD  n26 n180 DP_OP_94J1_122_9915_n238 XNOR2xp5_ASAP7_75t_R
XU278 VSS VDD  n182 n146 n180 XOR2xp5_ASAP7_75t_R
XU279 VSS VDD  in[41] n183 n182 XNOR2xp5_ASAP7_75t_R
XU280 VSS VDD  DP_OP_94J1_122_9915_n291 DP_OP_94J1_122_9915_n289 n184 XNOR2xp5_ASAP7_75t_R
XU281 VSS VDD  n97 DP_OP_94J1_122_9915_n100 n185 XNOR2xp5_ASAP7_75t_R
XU282 VSS VDD  DP_OP_94J1_122_9915_n274 DP_OP_94J1_122_9915_n276 DP_OP_94J1_122_9915_n238 DP_OP_94J1_122_9915_n226 MAJIxp5_ASAP7_75t_R
XU283 VSS VDD  n25 n98 n187 XOR2xp5_ASAP7_75t_R
XU284 VSS VDD  n188 n213 out[2] XNOR2xp5_ASAP7_75t_R
XU285 VSS VDD  n133 n211 n209 n188 MAJIxp5_ASAP7_75t_R
XU286 VSS VDD  DP_OP_94J1_122_9915_n146 DP_OP_94J1_122_9915_n142 DP_OP_94J1_122_9915_n148 DP_OP_94J1_122_9915_n117 MAJIxp5_ASAP7_75t_R
XU287 VSS VDD  DP_OP_94J1_122_9915_n62 n189 DP_OP_94J1_122_9915_n57 XOR2xp5_ASAP7_75t_R
XU288 VSS VDD  DP_OP_94J1_122_9915_n93 DP_OP_94J1_122_9915_n64 n189 XNOR2xp5_ASAP7_75t_R
XU289 VSS VDD  DP_OP_94J1_122_9915_n47 DP_OP_94J1_122_9915_n61 n196 NAND2xp33_ASAP7_75t_R
XU290 VSS VDD  in[110] in[118] in[42] DP_OP_94J1_122_9915_n203 MAJIxp5_ASAP7_75t_R
XU291 VSS VDD  in[110] n190 DP_OP_94J1_122_9915_n204 XNOR2xp5_ASAP7_75t_R
XU292 VSS VDD  in[2] n191 DP_OP_94J1_122_9915_n212 XNOR2xp5_ASAP7_75t_R
XU293 VSS VDD  in[45] in[61] in[53] DP_OP_94J1_122_9915_n265 MAJIxp5_ASAP7_75t_R
XU294 VSS VDD  in[45] n192 DP_OP_94J1_122_9915_n266 XNOR2xp5_ASAP7_75t_R
XU295 VSS VDD  DP_OP_94J1_122_9915_n277 DP_OP_94J1_122_9915_n275 DP_OP_94J1_122_9915_n273 n211 MAJIxp5_ASAP7_75t_R
XU296 VSS VDD  DP_OP_94J1_122_9915_n47 DP_OP_94J1_122_9915_n61 n198 OR2x2_ASAP7_75t_R
XU297 VSS VDD  in[24] in[16] in[8] DP_OP_94J1_122_9915_n281 MAJIxp5_ASAP7_75t_R
XU298 VSS VDD  in[24] n199 DP_OP_94J1_122_9915_n282 XNOR2xp5_ASAP7_75t_R
XU299 VSS VDD  in[47] in[55] in[115] DP_OP_94J1_122_9915_n151 MAJIxp5_ASAP7_75t_R
XU300 VSS VDD  DP_OP_94J1_122_9915_n244 n31 n202 XNOR2xp5_ASAP7_75t_R
XU301 VSS VDD  in[105] in[73] in[33] DP_OP_94J1_122_9915_n251 MAJIxp5_ASAP7_75t_R
XU302 VSS VDD  in[105] n203 DP_OP_94J1_122_9915_n252 XNOR2xp5_ASAP7_75t_R
XU303 VSS VDD  in[117] in[1] in[81] DP_OP_94J1_122_9915_n259 MAJIxp5_ASAP7_75t_R
XU304 VSS VDD  in[39] in[31] n205 XOR2x1_ASAP7_75t_R
XU305 VSS VDD  in[113] in[25] in[97] DP_OP_94J1_122_9915_n253 MAJIxp5_ASAP7_75t_R
XU306 VSS VDD  in[113] n206 DP_OP_94J1_122_9915_n254 XNOR2xp5_ASAP7_75t_R
XU307 VSS VDD  in[58] in[66] in[90] DP_OP_94J1_122_9915_n199 MAJIxp5_ASAP7_75t_R
XU308 VSS VDD  in[58] n207 DP_OP_94J1_122_9915_n200 XNOR2xp5_ASAP7_75t_R
XU309 VSS VDD  DP_OP_94J1_122_9915_n277 DP_OP_94J1_122_9915_n275 A3  n208 HAxp5_ASAP7_75t_R
XU310 VSS VDD  DP_OP_94J1_122_9915_n273 n208 A4  out[0] HAxp5_ASAP7_75t_R
XU311 VSS VDD  n209 DP_OP_94J1_122_9915_n222 A5  n210 HAxp5_ASAP7_75t_R
XU312 VSS VDD  n210 n211 A6  out[1] HAxp5_ASAP7_75t_R
XU313 VSS VDD  DP_OP_94J1_122_9915_n161 n212 n213 XOR2xp5_ASAP7_75t_R
XU314 VSS VDD  n73 n214 A7  out[3] HAxp5_ASAP7_75t_R
XU315 VSS VDD  n218 n143 A8  out[5] HAxp5_ASAP7_75t_R
XU316 VSS VDD  in[23] in[39] in[31] n222 MAJIxp5_ASAP7_75t_R
XU317 VSS VDD  n222 n221 DP_OP_94J1_122_9915_n83 NOR2xp33_ASAP7_75t_R
XU318 VSS VDD  n222 n221 DP_OP_94J1_122_9915_n84 XOR2xp5_ASAP7_75t_R
XU319 VSS VDD  DP_OP_94J1_122_9915_n51 DP_OP_94J1_122_9915_n36 INVx1_ASAP7_75t_R
XU320 VSS VDD  in[57] in[49] in[41] DP_OP_94J1_122_9915_n249 MAJIxp5_ASAP7_75t_R
XU321 VSS VDD  DP_OP_94J1_122_9915_n37 n154 A9  n223 HAxp5_ASAP7_75t_R
.ENDS


