.TITLE DIC_Final

***-----------------------***
***        setting        ***
***-----------------------***

.protect
.include '../08_TECH/LIB/7nm_TT.pm'
.include '../08_TECH/LIB/16mos.pm'
.include '../08_TECH/LIB/asap7sc7p5t_SIMPLE_RVT.sp' 
.include '../08_TECH/LIB/asap7sc7p5t_SEQ_RVT.sp'    
.include '../08_TECH/LIB/asap7sc7p5t_INVBUF_RVT.sp' 
.include '../08_TECH/LIB/asap7sc7p5t_AO_RVT.sp'     
.include '../08_TECH/LIB/asap7sc7p5t_OA_RVT.sp'     
.unprotect

.VEC "mul.vec" 

*** Voltage: 0.7V ***
.PARAM supply=0.7v

*** Temperature: 25C ***
.TEMP 25

***********************************
* Transition Analysis             *
***********************************
.TRAN 1ps 20ns 

***********************************
* HSPICE Options                  *
***********************************
.OPTION POST PROBE
.OPTION NOMOD BRIEF MEASDGT=7 
.OPTION CAPTAB NOTOP AUTOSTOP

***********************************
* Output Signals                  *
***********************************
.probe tran v(*) i(*)


***********************************
* Define Global Nets              *
***********************************
.GLOBAL VDD GND BL BLB

***********************************
* Voltage Sources                 *
***********************************
vdd     VDD   0  DC supply
vss     VSS   0  DC 0
vbl     BL    0   DC supply/2
vblb    BLB   0   DC supply/2

***********************************
* Measurement Commands            *
***********************************
.meas pwr avg POWER



***-----------------------***
***        circuit        ***
***-----------------------***


* // Xbuf Input In_bar INV
* // ADD INPUT BUFFER
* // WEIGHT IS INITIALIZE IN THE SRAM
* // SO CIM OPERATION IS READ THE WEIGHT AND THEN DO DOT PRODUCT 
* XI11 I111 I111_inv INV
* XI12 I112 I112_inv INV
* XI13 I113 I113_inv INV
* XI14 I114 I114_inv INV
* XI15 I121 I121_inv INV
* XI16 I122 I122_inv INV
* XI17 I123 I123_inv INV
* XI18 I124 I124_inv INV
* XI19 I131 I131_inv INV
* XI20 I132 I132_inv INV
* XI21 I133 I133_inv INV
* XI22 I134 I134_inv INV
* XI23 I141 I141_inv INV
* XI24 I142 I142_inv INV
* XI25 I143 I143_inv INV
* XI26 I144 I144_inv INV
* XI27 I151 I151_inv INV
* XI28 I152 I152_inv INV
* XI29 I153 I153_inv INV
* XI30 I154 I154_inv INV
* XI31 I161 I161_inv INV
* XI32 I162 I162_inv INV
* XI33 I163 I163_inv INV
* XI34 I164 I164_inv INV
* XI35 I171 I171_inv INV
* XI36 I172 I172_inv INV
* XI37 I173 I173_inv INV
* XI38 I174 I174_inv INV
* XI39 I181 I181_inv INV
* XI40 I182 I182_inv INV
* XI41 I183 I183_inv INV
* XI42 I184 I184_inv INV
* XI43 I191 I191_inv INV
* XI44 I192 I192_inv INV
* XI45 I193 I193_inv INV
* XI46 I194 I194_inv INV
* XI47 I1101 I1101_inv INV
* XI48 I1102 I1102_inv INV
* XI49 I1103 I1103_inv INV
* XI50 I1104 I1104_inv INV
* XI51 I1111 I1111_inv INV
* XI52 I1112 I1112_inv INV
* XI53 I1113 I1113_inv INV
* XI54 I1114 I1114_inv INV
* XI55 I1121 I1121_inv INV
* XI56 I1122 I1122_inv INV
* XI57 I1123 I1123_inv INV
* XI58 I1124 I1124_inv INV
* XI59 I1131 I1131_inv INV
* XI60 I1132 I1132_inv INV
* XI61 I1133 I1133_inv INV
* XI62 I1134 I1134_inv INV
* XI63 I1141 I1141_inv INV
* XI64 I1142 I1142_inv INV
* XI65 I1143 I1143_inv INV
* XI66 I1144 I1144_inv INV
* XI67 I1151 I1151_inv INV
* XI68 I1152 I1152_inv INV
* XI69 I1153 I1153_inv INV
* XI70 I1154 I1154_inv INV
* XI71 I1161 I1161_inv INV
* XI72 I1162 I1162_inv INV
* XI73 I1163 I1163_inv INV
* XI74 I1164 I1164_inv INV
* XI75 I1171 I1171_inv INV
* XI76 I1172 I1172_inv INV
* XI77 I1173 I1173_inv INV
* XI78 I1174 I1174_inv INV
* XI79 I1181 I1181_inv INV
* XI80 I1182 I1182_inv INV
* XI81 I1183 I1183_inv INV
* XI82 I1184 I1184_inv INV
* XI83 I1191 I1191_inv INV
* XI84 I1192 I1192_inv INV
* XI85 I1193 I1193_inv INV
* XI86 I1194 I1194_inv INV
* XI87 I1201 I1201_inv INV
* XI88 I1202 I1202_inv INV
* XI89 I1203 I1203_inv INV
* XI90 I1204 I1204_inv INV
* XI91 I1211 I1211_inv INV
* XI92 I1212 I1212_inv INV
* XI93 I1213 I1213_inv INV
* XI94 I1214 I1214_inv INV
* XI95 I1221 I1221_inv INV
* XI96 I1222 I1222_inv INV
* XI97 I1223 I1223_inv INV
* XI98 I1224 I1224_inv INV
* XI99 I1231 I1231_inv INV
* XI100 I1232 I1232_inv INV
* XI101 I1233 I1233_inv INV
* XI102 I1234 I1234_inv INV
* XI103 I1241 I1241_inv INV
* XI104 I1242 I1242_inv INV
* XI105 I1243 I1243_inv INV
* XI106 I1244 I1244_inv INV
* XI107 I1251 I1251_inv INV
* XI108 I1252 I1252_inv INV
* XI109 I1253 I1253_inv INV
* XI110 I1254 I1254_inv INV
* XI111 I1261 I1261_inv INV
* XI112 I1262 I1262_inv INV
* XI113 I1263 I1263_inv INV
* XI114 I1264 I1264_inv INV
* XI115 I1271 I1271_inv INV
* XI116 I1272 I1272_inv INV
* XI117 I1273 I1273_inv INV
* XI118 I1274 I1274_inv INV
* XI119 I1281 I1281_inv INV
* XI120 I1282 I1282_inv INV
* XI121 I1283 I1283_inv INV
* XI122 I1284 I1284_inv INV
* XI123 I1291 I1291_inv INV
* XI124 I1292 I1292_inv INV
* XI125 I1293 I1293_inv INV
* XI126 I1294 I1294_inv INV
* XI127 I1301 I1301_inv INV
* XI128 I1302 I1302_inv INV
* XI129 I1303 I1303_inv INV
* XI130 I1304 I1304_inv INV
* XI131 I1311 I1311_inv INV
* XI132 I1312 I1312_inv INV
* XI133 I1313 I1313_inv INV
* XI134 I1314 I1314_inv INV
* XI135 I1321 I1321_inv INV
* XI136 I1322 I1322_inv INV
* XI137 I1323 I1323_inv INV
* XI138 I1324 I1324_inv INV
* XI139 I211 I211_inv INV
* XI140 I212 I212_inv INV
* XI141 I213 I213_inv INV
* XI142 I214 I214_inv INV
* XI143 I221 I221_inv INV
* XI144 I222 I222_inv INV
* XI145 I223 I223_inv INV
* XI146 I224 I224_inv INV
* XI147 I231 I231_inv INV
* XI148 I232 I232_inv INV
* XI149 I233 I233_inv INV
* XI150 I234 I234_inv INV
* XI151 I241 I241_inv INV
* XI152 I242 I242_inv INV
* XI153 I243 I243_inv INV
* XI154 I244 I244_inv INV
* XI155 I251 I251_inv INV
* XI156 I252 I252_inv INV
* XI157 I253 I253_inv INV
* XI158 I254 I254_inv INV
* XI159 I261 I261_inv INV
* XI160 I262 I262_inv INV
* XI161 I263 I263_inv INV
* XI162 I264 I264_inv INV
* XI163 I271 I271_inv INV
* XI164 I272 I272_inv INV
* XI165 I273 I273_inv INV
* XI166 I274 I274_inv INV
* XI167 I281 I281_inv INV
* XI168 I282 I282_inv INV
* XI169 I283 I283_inv INV
* XI170 I284 I284_inv INV
* XI171 I291 I291_inv INV
* XI172 I292 I292_inv INV
* XI173 I293 I293_inv INV
* XI174 I294 I294_inv INV
* XI175 I2101 I2101_inv INV
* XI176 I2102 I2102_inv INV
* XI177 I2103 I2103_inv INV
* XI178 I2104 I2104_inv INV
* XI179 I2111 I2111_inv INV
* XI180 I2112 I2112_inv INV
* XI181 I2113 I2113_inv INV
* XI182 I2114 I2114_inv INV
* XI183 I2121 I2121_inv INV
* XI184 I2122 I2122_inv INV
* XI185 I2123 I2123_inv INV
* XI186 I2124 I2124_inv INV
* XI187 I2131 I2131_inv INV
* XI188 I2132 I2132_inv INV
* XI189 I2133 I2133_inv INV
* XI190 I2134 I2134_inv INV
* XI191 I2141 I2141_inv INV
* XI192 I2142 I2142_inv INV
* XI193 I2143 I2143_inv INV
* XI194 I2144 I2144_inv INV
* XI195 I2151 I2151_inv INV
* XI196 I2152 I2152_inv INV
* XI197 I2153 I2153_inv INV
* XI198 I2154 I2154_inv INV
* XI199 I2161 I2161_inv INV
* XI200 I2162 I2162_inv INV
* XI201 I2163 I2163_inv INV
* XI202 I2164 I2164_inv INV
* XI203 I2171 I2171_inv INV
* XI204 I2172 I2172_inv INV
* XI205 I2173 I2173_inv INV
* XI206 I2174 I2174_inv INV
* XI207 I2181 I2181_inv INV
* XI208 I2182 I2182_inv INV
* XI209 I2183 I2183_inv INV
* XI210 I2184 I2184_inv INV
* XI211 I2191 I2191_inv INV
* XI212 I2192 I2192_inv INV
* XI213 I2193 I2193_inv INV
* XI214 I2194 I2194_inv INV
* XI215 I2201 I2201_inv INV
* XI216 I2202 I2202_inv INV
* XI217 I2203 I2203_inv INV
* XI218 I2204 I2204_inv INV
* XI219 I2211 I2211_inv INV
* XI220 I2212 I2212_inv INV
* XI221 I2213 I2213_inv INV
* XI222 I2214 I2214_inv INV
* XI223 I2221 I2221_inv INV
* XI224 I2222 I2222_inv INV
* XI225 I2223 I2223_inv INV
* XI226 I2224 I2224_inv INV
* XI227 I2231 I2231_inv INV
* XI228 I2232 I2232_inv INV
* XI229 I2233 I2233_inv INV
* XI230 I2234 I2234_inv INV
* XI231 I2241 I2241_inv INV
* XI232 I2242 I2242_inv INV
* XI233 I2243 I2243_inv INV
* XI234 I2244 I2244_inv INV
* XI235 I2251 I2251_inv INV
* XI236 I2252 I2252_inv INV
* XI237 I2253 I2253_inv INV
* XI238 I2254 I2254_inv INV
* XI239 I2261 I2261_inv INV
* XI240 I2262 I2262_inv INV
* XI241 I2263 I2263_inv INV
* XI242 I2264 I2264_inv INV
* XI243 I2271 I2271_inv INV
* XI244 I2272 I2272_inv INV
* XI245 I2273 I2273_inv INV
* XI246 I2274 I2274_inv INV
* XI247 I2281 I2281_inv INV
* XI248 I2282 I2282_inv INV
* XI249 I2283 I2283_inv INV
* XI250 I2284 I2284_inv INV
* XI251 I2291 I2291_inv INV
* XI252 I2292 I2292_inv INV
* XI253 I2293 I2293_inv INV
* XI254 I2294 I2294_inv INV
* XI255 I2301 I2301_inv INV
* XI256 I2302 I2302_inv INV
* XI257 I2303 I2303_inv INV
* XI258 I2304 I2304_inv INV
* XI259 I2311 I2311_inv INV
* XI260 I2312 I2312_inv INV
* XI261 I2313 I2313_inv INV
* XI262 I2314 I2314_inv INV
* XI263 I2321 I2321_inv INV
* XI264 I2322 I2322_inv INV
* XI265 I2323 I2323_inv INV
* XI266 I2324 I2324_inv INV
* XI267 I311 I311_inv INV
* XI268 I312 I312_inv INV
* XI269 I313 I313_inv INV
* XI270 I314 I314_inv INV
* XI271 I321 I321_inv INV
* XI272 I322 I322_inv INV
* XI273 I323 I323_inv INV
* XI274 I324 I324_inv INV
* XI275 I331 I331_inv INV
* XI276 I332 I332_inv INV
* XI277 I333 I333_inv INV
* XI278 I334 I334_inv INV
* XI279 I341 I341_inv INV
* XI280 I342 I342_inv INV
* XI281 I343 I343_inv INV
* XI282 I344 I344_inv INV
* XI283 I351 I351_inv INV
* XI284 I352 I352_inv INV
* XI285 I353 I353_inv INV
* XI286 I354 I354_inv INV
* XI287 I361 I361_inv INV
* XI288 I362 I362_inv INV
* XI289 I363 I363_inv INV
* XI290 I364 I364_inv INV
* XI291 I371 I371_inv INV
* XI292 I372 I372_inv INV
* XI293 I373 I373_inv INV
* XI294 I374 I374_inv INV
* XI295 I381 I381_inv INV
* XI296 I382 I382_inv INV
* XI297 I383 I383_inv INV
* XI298 I384 I384_inv INV
* XI299 I391 I391_inv INV
* XI300 I392 I392_inv INV
* XI301 I393 I393_inv INV
* XI302 I394 I394_inv INV
* XI303 I3101 I3101_inv INV
* XI304 I3102 I3102_inv INV
* XI305 I3103 I3103_inv INV
* XI306 I3104 I3104_inv INV
* XI307 I3111 I3111_inv INV
* XI308 I3112 I3112_inv INV
* XI309 I3113 I3113_inv INV
* XI310 I3114 I3114_inv INV
* XI311 I3121 I3121_inv INV
* XI312 I3122 I3122_inv INV
* XI313 I3123 I3123_inv INV
* XI314 I3124 I3124_inv INV
* XI315 I3131 I3131_inv INV
* XI316 I3132 I3132_inv INV
* XI317 I3133 I3133_inv INV
* XI318 I3134 I3134_inv INV
* XI319 I3141 I3141_inv INV
* XI320 I3142 I3142_inv INV
* XI321 I3143 I3143_inv INV
* XI322 I3144 I3144_inv INV
* XI323 I3151 I3151_inv INV
* XI324 I3152 I3152_inv INV
* XI325 I3153 I3153_inv INV
* XI326 I3154 I3154_inv INV
* XI327 I3161 I3161_inv INV
* XI328 I3162 I3162_inv INV
* XI329 I3163 I3163_inv INV
* XI330 I3164 I3164_inv INV
* XI331 I3171 I3171_inv INV
* XI332 I3172 I3172_inv INV
* XI333 I3173 I3173_inv INV
* XI334 I3174 I3174_inv INV
* XI335 I3181 I3181_inv INV
* XI336 I3182 I3182_inv INV
* XI337 I3183 I3183_inv INV
* XI338 I3184 I3184_inv INV
* XI339 I3191 I3191_inv INV
* XI340 I3192 I3192_inv INV
* XI341 I3193 I3193_inv INV
* XI342 I3194 I3194_inv INV
* XI343 I3201 I3201_inv INV
* XI344 I3202 I3202_inv INV
* XI345 I3203 I3203_inv INV
* XI346 I3204 I3204_inv INV
* XI347 I3211 I3211_inv INV
* XI348 I3212 I3212_inv INV
* XI349 I3213 I3213_inv INV
* XI350 I3214 I3214_inv INV
* XI351 I3221 I3221_inv INV
* XI352 I3222 I3222_inv INV
* XI353 I3223 I3223_inv INV
* XI354 I3224 I3224_inv INV
* XI355 I3231 I3231_inv INV
* XI356 I3232 I3232_inv INV
* XI357 I3233 I3233_inv INV
* XI358 I3234 I3234_inv INV
* XI359 I3241 I3241_inv INV
* XI360 I3242 I3242_inv INV
* XI361 I3243 I3243_inv INV
* XI362 I3244 I3244_inv INV
* XI363 I3251 I3251_inv INV
* XI364 I3252 I3252_inv INV
* XI365 I3253 I3253_inv INV
* XI366 I3254 I3254_inv INV
* XI367 I3261 I3261_inv INV
* XI368 I3262 I3262_inv INV
* XI369 I3263 I3263_inv INV
* XI370 I3264 I3264_inv INV
* XI371 I3271 I3271_inv INV
* XI372 I3272 I3272_inv INV
* XI373 I3273 I3273_inv INV
* XI374 I3274 I3274_inv INV
* XI375 I3281 I3281_inv INV
* XI376 I3282 I3282_inv INV
* XI377 I3283 I3283_inv INV
* XI378 I3284 I3284_inv INV
* XI379 I3291 I3291_inv INV
* XI380 I3292 I3292_inv INV
* XI381 I3293 I3293_inv INV
* XI382 I3294 I3294_inv INV
* XI383 I3301 I3301_inv INV
* XI384 I3302 I3302_inv INV
* XI385 I3303 I3303_inv INV
* XI386 I3304 I3304_inv INV
* XI387 I3311 I3311_inv INV
* XI388 I3312 I3312_inv INV
* XI389 I3313 I3313_inv INV
* XI390 I3314 I3314_inv INV
* XI391 I3321 I3321_inv INV
* XI392 I3322 I3322_inv INV
* XI393 I3323 I3323_inv INV
* XI394 I3324 I3324_inv INV
* XI395 I411 I411_inv INV
* XI396 I412 I412_inv INV
* XI397 I413 I413_inv INV
* XI398 I414 I414_inv INV
* XI399 I421 I421_inv INV
* XI400 I422 I422_inv INV
* XI401 I423 I423_inv INV
* XI402 I424 I424_inv INV
* XI403 I431 I431_inv INV
* XI404 I432 I432_inv INV
* XI405 I433 I433_inv INV
* XI406 I434 I434_inv INV
* XI407 I441 I441_inv INV
* XI408 I442 I442_inv INV
* XI409 I443 I443_inv INV
* XI410 I444 I444_inv INV
* XI411 I451 I451_inv INV
* XI412 I452 I452_inv INV
* XI413 I453 I453_inv INV
* XI414 I454 I454_inv INV
* XI415 I461 I461_inv INV
* XI416 I462 I462_inv INV
* XI417 I463 I463_inv INV
* XI418 I464 I464_inv INV
* XI419 I471 I471_inv INV
* XI420 I472 I472_inv INV
* XI421 I473 I473_inv INV
* XI422 I474 I474_inv INV
* XI423 I481 I481_inv INV
* XI424 I482 I482_inv INV
* XI425 I483 I483_inv INV
* XI426 I484 I484_inv INV
* XI427 I491 I491_inv INV
* XI428 I492 I492_inv INV
* XI429 I493 I493_inv INV
* XI430 I494 I494_inv INV
* XI431 I4101 I4101_inv INV
* XI432 I4102 I4102_inv INV
* XI433 I4103 I4103_inv INV
* XI434 I4104 I4104_inv INV
* XI435 I4111 I4111_inv INV
* XI436 I4112 I4112_inv INV
* XI437 I4113 I4113_inv INV
* XI438 I4114 I4114_inv INV
* XI439 I4121 I4121_inv INV
* XI440 I4122 I4122_inv INV
* XI441 I4123 I4123_inv INV
* XI442 I4124 I4124_inv INV
* XI443 I4131 I4131_inv INV
* XI444 I4132 I4132_inv INV
* XI445 I4133 I4133_inv INV
* XI446 I4134 I4134_inv INV
* XI447 I4141 I4141_inv INV
* XI448 I4142 I4142_inv INV
* XI449 I4143 I4143_inv INV
* XI450 I4144 I4144_inv INV
* XI451 I4151 I4151_inv INV
* XI452 I4152 I4152_inv INV
* XI453 I4153 I4153_inv INV
* XI454 I4154 I4154_inv INV
* XI455 I4161 I4161_inv INV
* XI456 I4162 I4162_inv INV
* XI457 I4163 I4163_inv INV
* XI458 I4164 I4164_inv INV
* XI459 I4171 I4171_inv INV
* XI460 I4172 I4172_inv INV
* XI461 I4173 I4173_inv INV
* XI462 I4174 I4174_inv INV
* XI463 I4181 I4181_inv INV
* XI464 I4182 I4182_inv INV
* XI465 I4183 I4183_inv INV
* XI466 I4184 I4184_inv INV
* XI467 I4191 I4191_inv INV
* XI468 I4192 I4192_inv INV
* XI469 I4193 I4193_inv INV
* XI470 I4194 I4194_inv INV
* XI471 I4201 I4201_inv INV
* XI472 I4202 I4202_inv INV
* XI473 I4203 I4203_inv INV
* XI474 I4204 I4204_inv INV
* XI475 I4211 I4211_inv INV
* XI476 I4212 I4212_inv INV
* XI477 I4213 I4213_inv INV
* XI478 I4214 I4214_inv INV
* XI479 I4221 I4221_inv INV
* XI480 I4222 I4222_inv INV
* XI481 I4223 I4223_inv INV
* XI482 I4224 I4224_inv INV
* XI483 I4231 I4231_inv INV
* XI484 I4232 I4232_inv INV
* XI485 I4233 I4233_inv INV
* XI486 I4234 I4234_inv INV
* XI487 I4241 I4241_inv INV
* XI488 I4242 I4242_inv INV
* XI489 I4243 I4243_inv INV
* XI490 I4244 I4244_inv INV
* XI491 I4251 I4251_inv INV
* XI492 I4252 I4252_inv INV
* XI493 I4253 I4253_inv INV
* XI494 I4254 I4254_inv INV
* XI495 I4261 I4261_inv INV
* XI496 I4262 I4262_inv INV
* XI497 I4263 I4263_inv INV
* XI498 I4264 I4264_inv INV
* XI499 I4271 I4271_inv INV
* XI500 I4272 I4272_inv INV
* XI501 I4273 I4273_inv INV
* XI502 I4274 I4274_inv INV
* XI503 I4281 I4281_inv INV
* XI504 I4282 I4282_inv INV
* XI505 I4283 I4283_inv INV
* XI506 I4284 I4284_inv INV
* XI507 I4291 I4291_inv INV
* XI508 I4292 I4292_inv INV
* XI509 I4293 I4293_inv INV
* XI510 I4294 I4294_inv INV
* XI511 I4301 I4301_inv INV
* XI512 I4302 I4302_inv INV
* XI513 I4303 I4303_inv INV
* XI514 I4304 I4304_inv INV
* XI515 I4311 I4311_inv INV
* XI516 I4312 I4312_inv INV
* XI517 I4313 I4313_inv INV
* XI518 I4314 I4314_inv INV
* XI519 I4321 I4321_inv INV
* XI520 I4322 I4322_inv INV
* XI521 I4323 I4323_inv INV
* XI522 I4324 I4324_inv INV

XI11 I111 I111_buf INV
XB11 I111_buf I111_inv Buffer
XI12 I112 I112_buf INV
XB12 I112_buf I112_inv Buffer
XI13 I113 I113_buf INV
XB13 I113_buf I113_inv Buffer
XI14 I114 I114_buf INV
XB14 I114_buf I114_inv Buffer
XI15 I121 I121_buf INV
XB15 I121_buf I121_inv Buffer
XI16 I122 I122_buf INV
XB16 I122_buf I122_inv Buffer
XI17 I123 I123_buf INV
XB17 I123_buf I123_inv Buffer
XI18 I124 I124_buf INV
XB18 I124_buf I124_inv Buffer
XI19 I131 I131_buf INV
XB19 I131_buf I131_inv Buffer
XI20 I132 I132_buf INV
XB20 I132_buf I132_inv Buffer
XI21 I133 I133_buf INV
XB21 I133_buf I133_inv Buffer
XI22 I134 I134_buf INV
XB22 I134_buf I134_inv Buffer
XI23 I141 I141_buf INV
XB23 I141_buf I141_inv Buffer
XI24 I142 I142_buf INV
XB24 I142_buf I142_inv Buffer
XI25 I143 I143_buf INV
XB25 I143_buf I143_inv Buffer
XI26 I144 I144_buf INV
XB26 I144_buf I144_inv Buffer
XI27 I151 I151_buf INV
XB27 I151_buf I151_inv Buffer
XI28 I152 I152_buf INV
XB28 I152_buf I152_inv Buffer
XI29 I153 I153_buf INV
XB29 I153_buf I153_inv Buffer
XI30 I154 I154_buf INV
XB30 I154_buf I154_inv Buffer
XI31 I161 I161_buf INV
XB31 I161_buf I161_inv Buffer
XI32 I162 I162_buf INV
XB32 I162_buf I162_inv Buffer
XI33 I163 I163_buf INV
XB33 I163_buf I163_inv Buffer
XI34 I164 I164_buf INV
XB34 I164_buf I164_inv Buffer
XI35 I171 I171_buf INV
XB35 I171_buf I171_inv Buffer
XI36 I172 I172_buf INV
XB36 I172_buf I172_inv Buffer
XI37 I173 I173_buf INV
XB37 I173_buf I173_inv Buffer
XI38 I174 I174_buf INV
XB38 I174_buf I174_inv Buffer
XI39 I181 I181_buf INV
XB39 I181_buf I181_inv Buffer
XI40 I182 I182_buf INV
XB40 I182_buf I182_inv Buffer
XI41 I183 I183_buf INV
XB41 I183_buf I183_inv Buffer
XI42 I184 I184_buf INV
XB42 I184_buf I184_inv Buffer
XI43 I191 I191_buf INV
XB43 I191_buf I191_inv Buffer
XI44 I192 I192_buf INV
XB44 I192_buf I192_inv Buffer
XI45 I193 I193_buf INV
XB45 I193_buf I193_inv Buffer
XI46 I194 I194_buf INV
XB46 I194_buf I194_inv Buffer
XI47 I1101 I1101_buf INV
XB47 I1101_buf I1101_inv Buffer
XI48 I1102 I1102_buf INV
XB48 I1102_buf I1102_inv Buffer
XI49 I1103 I1103_buf INV
XB49 I1103_buf I1103_inv Buffer
XI50 I1104 I1104_buf INV
XB50 I1104_buf I1104_inv Buffer
XI51 I1111 I1111_buf INV
XB51 I1111_buf I1111_inv Buffer
XI52 I1112 I1112_buf INV
XB52 I1112_buf I1112_inv Buffer
XI53 I1113 I1113_buf INV
XB53 I1113_buf I1113_inv Buffer
XI54 I1114 I1114_buf INV
XB54 I1114_buf I1114_inv Buffer
XI55 I1121 I1121_buf INV
XB55 I1121_buf I1121_inv Buffer
XI56 I1122 I1122_buf INV
XB56 I1122_buf I1122_inv Buffer
XI57 I1123 I1123_buf INV
XB57 I1123_buf I1123_inv Buffer
XI58 I1124 I1124_buf INV
XB58 I1124_buf I1124_inv Buffer
XI59 I1131 I1131_buf INV
XB59 I1131_buf I1131_inv Buffer
XI60 I1132 I1132_buf INV
XB60 I1132_buf I1132_inv Buffer
XI61 I1133 I1133_buf INV
XB61 I1133_buf I1133_inv Buffer
XI62 I1134 I1134_buf INV
XB62 I1134_buf I1134_inv Buffer
XI63 I1141 I1141_buf INV
XB63 I1141_buf I1141_inv Buffer
XI64 I1142 I1142_buf INV
XB64 I1142_buf I1142_inv Buffer
XI65 I1143 I1143_buf INV
XB65 I1143_buf I1143_inv Buffer
XI66 I1144 I1144_buf INV
XB66 I1144_buf I1144_inv Buffer
XI67 I1151 I1151_buf INV
XB67 I1151_buf I1151_inv Buffer
XI68 I1152 I1152_buf INV
XB68 I1152_buf I1152_inv Buffer
XI69 I1153 I1153_buf INV
XB69 I1153_buf I1153_inv Buffer
XI70 I1154 I1154_buf INV
XB70 I1154_buf I1154_inv Buffer
XI71 I1161 I1161_buf INV
XB71 I1161_buf I1161_inv Buffer
XI72 I1162 I1162_buf INV
XB72 I1162_buf I1162_inv Buffer
XI73 I1163 I1163_buf INV
XB73 I1163_buf I1163_inv Buffer
XI74 I1164 I1164_buf INV
XB74 I1164_buf I1164_inv Buffer
XI75 I1171 I1171_buf INV
XB75 I1171_buf I1171_inv Buffer
XI76 I1172 I1172_buf INV
XB76 I1172_buf I1172_inv Buffer
XI77 I1173 I1173_buf INV
XB77 I1173_buf I1173_inv Buffer
XI78 I1174 I1174_buf INV
XB78 I1174_buf I1174_inv Buffer
XI79 I1181 I1181_buf INV
XB79 I1181_buf I1181_inv Buffer
XI80 I1182 I1182_buf INV
XB80 I1182_buf I1182_inv Buffer
XI81 I1183 I1183_buf INV
XB81 I1183_buf I1183_inv Buffer
XI82 I1184 I1184_buf INV
XB82 I1184_buf I1184_inv Buffer
XI83 I1191 I1191_buf INV
XB83 I1191_buf I1191_inv Buffer
XI84 I1192 I1192_buf INV
XB84 I1192_buf I1192_inv Buffer
XI85 I1193 I1193_buf INV
XB85 I1193_buf I1193_inv Buffer
XI86 I1194 I1194_buf INV
XB86 I1194_buf I1194_inv Buffer
XI87 I1201 I1201_buf INV
XB87 I1201_buf I1201_inv Buffer
XI88 I1202 I1202_buf INV
XB88 I1202_buf I1202_inv Buffer
XI89 I1203 I1203_buf INV
XB89 I1203_buf I1203_inv Buffer
XI90 I1204 I1204_buf INV
XB90 I1204_buf I1204_inv Buffer
XI91 I1211 I1211_buf INV
XB91 I1211_buf I1211_inv Buffer
XI92 I1212 I1212_buf INV
XB92 I1212_buf I1212_inv Buffer
XI93 I1213 I1213_buf INV
XB93 I1213_buf I1213_inv Buffer
XI94 I1214 I1214_buf INV
XB94 I1214_buf I1214_inv Buffer
XI95 I1221 I1221_buf INV
XB95 I1221_buf I1221_inv Buffer
XI96 I1222 I1222_buf INV
XB96 I1222_buf I1222_inv Buffer
XI97 I1223 I1223_buf INV
XB97 I1223_buf I1223_inv Buffer
XI98 I1224 I1224_buf INV
XB98 I1224_buf I1224_inv Buffer
XI99 I1231 I1231_buf INV
XB99 I1231_buf I1231_inv Buffer
XI100 I1232 I1232_buf INV
XB100 I1232_buf I1232_inv Buffer
XI101 I1233 I1233_buf INV
XB101 I1233_buf I1233_inv Buffer
XI102 I1234 I1234_buf INV
XB102 I1234_buf I1234_inv Buffer
XI103 I1241 I1241_buf INV
XB103 I1241_buf I1241_inv Buffer
XI104 I1242 I1242_buf INV
XB104 I1242_buf I1242_inv Buffer
XI105 I1243 I1243_buf INV
XB105 I1243_buf I1243_inv Buffer
XI106 I1244 I1244_buf INV
XB106 I1244_buf I1244_inv Buffer
XI107 I1251 I1251_buf INV
XB107 I1251_buf I1251_inv Buffer
XI108 I1252 I1252_buf INV
XB108 I1252_buf I1252_inv Buffer
XI109 I1253 I1253_buf INV
XB109 I1253_buf I1253_inv Buffer
XI110 I1254 I1254_buf INV
XB110 I1254_buf I1254_inv Buffer
XI111 I1261 I1261_buf INV
XB111 I1261_buf I1261_inv Buffer
XI112 I1262 I1262_buf INV
XB112 I1262_buf I1262_inv Buffer
XI113 I1263 I1263_buf INV
XB113 I1263_buf I1263_inv Buffer
XI114 I1264 I1264_buf INV
XB114 I1264_buf I1264_inv Buffer
XI115 I1271 I1271_buf INV
XB115 I1271_buf I1271_inv Buffer
XI116 I1272 I1272_buf INV
XB116 I1272_buf I1272_inv Buffer
XI117 I1273 I1273_buf INV
XB117 I1273_buf I1273_inv Buffer
XI118 I1274 I1274_buf INV
XB118 I1274_buf I1274_inv Buffer
XI119 I1281 I1281_buf INV
XB119 I1281_buf I1281_inv Buffer
XI120 I1282 I1282_buf INV
XB120 I1282_buf I1282_inv Buffer
XI121 I1283 I1283_buf INV
XB121 I1283_buf I1283_inv Buffer
XI122 I1284 I1284_buf INV
XB122 I1284_buf I1284_inv Buffer
XI123 I1291 I1291_buf INV
XB123 I1291_buf I1291_inv Buffer
XI124 I1292 I1292_buf INV
XB124 I1292_buf I1292_inv Buffer
XI125 I1293 I1293_buf INV
XB125 I1293_buf I1293_inv Buffer
XI126 I1294 I1294_buf INV
XB126 I1294_buf I1294_inv Buffer
XI127 I1301 I1301_buf INV
XB127 I1301_buf I1301_inv Buffer
XI128 I1302 I1302_buf INV
XB128 I1302_buf I1302_inv Buffer
XI129 I1303 I1303_buf INV
XB129 I1303_buf I1303_inv Buffer
XI130 I1304 I1304_buf INV
XB130 I1304_buf I1304_inv Buffer
XI131 I1311 I1311_buf INV
XB131 I1311_buf I1311_inv Buffer
XI132 I1312 I1312_buf INV
XB132 I1312_buf I1312_inv Buffer
XI133 I1313 I1313_buf INV
XB133 I1313_buf I1313_inv Buffer
XI134 I1314 I1314_buf INV
XB134 I1314_buf I1314_inv Buffer
XI135 I1321 I1321_buf INV
XB135 I1321_buf I1321_inv Buffer
XI136 I1322 I1322_buf INV
XB136 I1322_buf I1322_inv Buffer
XI137 I1323 I1323_buf INV
XB137 I1323_buf I1323_inv Buffer
XI138 I1324 I1324_buf INV
XB138 I1324_buf I1324_inv Buffer
XI139 I211 I211_buf INV
XB139 I211_buf I211_inv Buffer
XI140 I212 I212_buf INV
XB140 I212_buf I212_inv Buffer
XI141 I213 I213_buf INV
XB141 I213_buf I213_inv Buffer
XI142 I214 I214_buf INV
XB142 I214_buf I214_inv Buffer
XI143 I221 I221_buf INV
XB143 I221_buf I221_inv Buffer
XI144 I222 I222_buf INV
XB144 I222_buf I222_inv Buffer
XI145 I223 I223_buf INV
XB145 I223_buf I223_inv Buffer
XI146 I224 I224_buf INV
XB146 I224_buf I224_inv Buffer
XI147 I231 I231_buf INV
XB147 I231_buf I231_inv Buffer
XI148 I232 I232_buf INV
XB148 I232_buf I232_inv Buffer
XI149 I233 I233_buf INV
XB149 I233_buf I233_inv Buffer
XI150 I234 I234_buf INV
XB150 I234_buf I234_inv Buffer
XI151 I241 I241_buf INV
XB151 I241_buf I241_inv Buffer
XI152 I242 I242_buf INV
XB152 I242_buf I242_inv Buffer
XI153 I243 I243_buf INV
XB153 I243_buf I243_inv Buffer
XI154 I244 I244_buf INV
XB154 I244_buf I244_inv Buffer
XI155 I251 I251_buf INV
XB155 I251_buf I251_inv Buffer
XI156 I252 I252_buf INV
XB156 I252_buf I252_inv Buffer
XI157 I253 I253_buf INV
XB157 I253_buf I253_inv Buffer
XI158 I254 I254_buf INV
XB158 I254_buf I254_inv Buffer
XI159 I261 I261_buf INV
XB159 I261_buf I261_inv Buffer
XI160 I262 I262_buf INV
XB160 I262_buf I262_inv Buffer
XI161 I263 I263_buf INV
XB161 I263_buf I263_inv Buffer
XI162 I264 I264_buf INV
XB162 I264_buf I264_inv Buffer
XI163 I271 I271_buf INV
XB163 I271_buf I271_inv Buffer
XI164 I272 I272_buf INV
XB164 I272_buf I272_inv Buffer
XI165 I273 I273_buf INV
XB165 I273_buf I273_inv Buffer
XI166 I274 I274_buf INV
XB166 I274_buf I274_inv Buffer
XI167 I281 I281_buf INV
XB167 I281_buf I281_inv Buffer
XI168 I282 I282_buf INV
XB168 I282_buf I282_inv Buffer
XI169 I283 I283_buf INV
XB169 I283_buf I283_inv Buffer
XI170 I284 I284_buf INV
XB170 I284_buf I284_inv Buffer
XI171 I291 I291_buf INV
XB171 I291_buf I291_inv Buffer
XI172 I292 I292_buf INV
XB172 I292_buf I292_inv Buffer
XI173 I293 I293_buf INV
XB173 I293_buf I293_inv Buffer
XI174 I294 I294_buf INV
XB174 I294_buf I294_inv Buffer
XI175 I2101 I2101_buf INV
XB175 I2101_buf I2101_inv Buffer
XI176 I2102 I2102_buf INV
XB176 I2102_buf I2102_inv Buffer
XI177 I2103 I2103_buf INV
XB177 I2103_buf I2103_inv Buffer
XI178 I2104 I2104_buf INV
XB178 I2104_buf I2104_inv Buffer
XI179 I2111 I2111_buf INV
XB179 I2111_buf I2111_inv Buffer
XI180 I2112 I2112_buf INV
XB180 I2112_buf I2112_inv Buffer
XI181 I2113 I2113_buf INV
XB181 I2113_buf I2113_inv Buffer
XI182 I2114 I2114_buf INV
XB182 I2114_buf I2114_inv Buffer
XI183 I2121 I2121_buf INV
XB183 I2121_buf I2121_inv Buffer
XI184 I2122 I2122_buf INV
XB184 I2122_buf I2122_inv Buffer
XI185 I2123 I2123_buf INV
XB185 I2123_buf I2123_inv Buffer
XI186 I2124 I2124_buf INV
XB186 I2124_buf I2124_inv Buffer
XI187 I2131 I2131_buf INV
XB187 I2131_buf I2131_inv Buffer
XI188 I2132 I2132_buf INV
XB188 I2132_buf I2132_inv Buffer
XI189 I2133 I2133_buf INV
XB189 I2133_buf I2133_inv Buffer
XI190 I2134 I2134_buf INV
XB190 I2134_buf I2134_inv Buffer
XI191 I2141 I2141_buf INV
XB191 I2141_buf I2141_inv Buffer
XI192 I2142 I2142_buf INV
XB192 I2142_buf I2142_inv Buffer
XI193 I2143 I2143_buf INV
XB193 I2143_buf I2143_inv Buffer
XI194 I2144 I2144_buf INV
XB194 I2144_buf I2144_inv Buffer
XI195 I2151 I2151_buf INV
XB195 I2151_buf I2151_inv Buffer
XI196 I2152 I2152_buf INV
XB196 I2152_buf I2152_inv Buffer
XI197 I2153 I2153_buf INV
XB197 I2153_buf I2153_inv Buffer
XI198 I2154 I2154_buf INV
XB198 I2154_buf I2154_inv Buffer
XI199 I2161 I2161_buf INV
XB199 I2161_buf I2161_inv Buffer
XI200 I2162 I2162_buf INV
XB200 I2162_buf I2162_inv Buffer
XI201 I2163 I2163_buf INV
XB201 I2163_buf I2163_inv Buffer
XI202 I2164 I2164_buf INV
XB202 I2164_buf I2164_inv Buffer
XI203 I2171 I2171_buf INV
XB203 I2171_buf I2171_inv Buffer
XI204 I2172 I2172_buf INV
XB204 I2172_buf I2172_inv Buffer
XI205 I2173 I2173_buf INV
XB205 I2173_buf I2173_inv Buffer
XI206 I2174 I2174_buf INV
XB206 I2174_buf I2174_inv Buffer
XI207 I2181 I2181_buf INV
XB207 I2181_buf I2181_inv Buffer
XI208 I2182 I2182_buf INV
XB208 I2182_buf I2182_inv Buffer
XI209 I2183 I2183_buf INV
XB209 I2183_buf I2183_inv Buffer
XI210 I2184 I2184_buf INV
XB210 I2184_buf I2184_inv Buffer
XI211 I2191 I2191_buf INV
XB211 I2191_buf I2191_inv Buffer
XI212 I2192 I2192_buf INV
XB212 I2192_buf I2192_inv Buffer
XI213 I2193 I2193_buf INV
XB213 I2193_buf I2193_inv Buffer
XI214 I2194 I2194_buf INV
XB214 I2194_buf I2194_inv Buffer
XI215 I2201 I2201_buf INV
XB215 I2201_buf I2201_inv Buffer
XI216 I2202 I2202_buf INV
XB216 I2202_buf I2202_inv Buffer
XI217 I2203 I2203_buf INV
XB217 I2203_buf I2203_inv Buffer
XI218 I2204 I2204_buf INV
XB218 I2204_buf I2204_inv Buffer
XI219 I2211 I2211_buf INV
XB219 I2211_buf I2211_inv Buffer
XI220 I2212 I2212_buf INV
XB220 I2212_buf I2212_inv Buffer
XI221 I2213 I2213_buf INV
XB221 I2213_buf I2213_inv Buffer
XI222 I2214 I2214_buf INV
XB222 I2214_buf I2214_inv Buffer
XI223 I2221 I2221_buf INV
XB223 I2221_buf I2221_inv Buffer
XI224 I2222 I2222_buf INV
XB224 I2222_buf I2222_inv Buffer
XI225 I2223 I2223_buf INV
XB225 I2223_buf I2223_inv Buffer
XI226 I2224 I2224_buf INV
XB226 I2224_buf I2224_inv Buffer
XI227 I2231 I2231_buf INV
XB227 I2231_buf I2231_inv Buffer
XI228 I2232 I2232_buf INV
XB228 I2232_buf I2232_inv Buffer
XI229 I2233 I2233_buf INV
XB229 I2233_buf I2233_inv Buffer
XI230 I2234 I2234_buf INV
XB230 I2234_buf I2234_inv Buffer
XI231 I2241 I2241_buf INV
XB231 I2241_buf I2241_inv Buffer
XI232 I2242 I2242_buf INV
XB232 I2242_buf I2242_inv Buffer
XI233 I2243 I2243_buf INV
XB233 I2243_buf I2243_inv Buffer
XI234 I2244 I2244_buf INV
XB234 I2244_buf I2244_inv Buffer
XI235 I2251 I2251_buf INV
XB235 I2251_buf I2251_inv Buffer
XI236 I2252 I2252_buf INV
XB236 I2252_buf I2252_inv Buffer
XI237 I2253 I2253_buf INV
XB237 I2253_buf I2253_inv Buffer
XI238 I2254 I2254_buf INV
XB238 I2254_buf I2254_inv Buffer
XI239 I2261 I2261_buf INV
XB239 I2261_buf I2261_inv Buffer
XI240 I2262 I2262_buf INV
XB240 I2262_buf I2262_inv Buffer
XI241 I2263 I2263_buf INV
XB241 I2263_buf I2263_inv Buffer
XI242 I2264 I2264_buf INV
XB242 I2264_buf I2264_inv Buffer
XI243 I2271 I2271_buf INV
XB243 I2271_buf I2271_inv Buffer
XI244 I2272 I2272_buf INV
XB244 I2272_buf I2272_inv Buffer
XI245 I2273 I2273_buf INV
XB245 I2273_buf I2273_inv Buffer
XI246 I2274 I2274_buf INV
XB246 I2274_buf I2274_inv Buffer
XI247 I2281 I2281_buf INV
XB247 I2281_buf I2281_inv Buffer
XI248 I2282 I2282_buf INV
XB248 I2282_buf I2282_inv Buffer
XI249 I2283 I2283_buf INV
XB249 I2283_buf I2283_inv Buffer
XI250 I2284 I2284_buf INV
XB250 I2284_buf I2284_inv Buffer
XI251 I2291 I2291_buf INV
XB251 I2291_buf I2291_inv Buffer
XI252 I2292 I2292_buf INV
XB252 I2292_buf I2292_inv Buffer
XI253 I2293 I2293_buf INV
XB253 I2293_buf I2293_inv Buffer
XI254 I2294 I2294_buf INV
XB254 I2294_buf I2294_inv Buffer
XI255 I2301 I2301_buf INV
XB255 I2301_buf I2301_inv Buffer
XI256 I2302 I2302_buf INV
XB256 I2302_buf I2302_inv Buffer
XI257 I2303 I2303_buf INV
XB257 I2303_buf I2303_inv Buffer
XI258 I2304 I2304_buf INV
XB258 I2304_buf I2304_inv Buffer
XI259 I2311 I2311_buf INV
XB259 I2311_buf I2311_inv Buffer
XI260 I2312 I2312_buf INV
XB260 I2312_buf I2312_inv Buffer
XI261 I2313 I2313_buf INV
XB261 I2313_buf I2313_inv Buffer
XI262 I2314 I2314_buf INV
XB262 I2314_buf I2314_inv Buffer
XI263 I2321 I2321_buf INV
XB263 I2321_buf I2321_inv Buffer
XI264 I2322 I2322_buf INV
XB264 I2322_buf I2322_inv Buffer
XI265 I2323 I2323_buf INV
XB265 I2323_buf I2323_inv Buffer
XI266 I2324 I2324_buf INV
XB266 I2324_buf I2324_inv Buffer
XI267 I311 I311_buf INV
XB267 I311_buf I311_inv Buffer
XI268 I312 I312_buf INV
XB268 I312_buf I312_inv Buffer
XI269 I313 I313_buf INV
XB269 I313_buf I313_inv Buffer
XI270 I314 I314_buf INV
XB270 I314_buf I314_inv Buffer
XI271 I321 I321_buf INV
XB271 I321_buf I321_inv Buffer
XI272 I322 I322_buf INV
XB272 I322_buf I322_inv Buffer
XI273 I323 I323_buf INV
XB273 I323_buf I323_inv Buffer
XI274 I324 I324_buf INV
XB274 I324_buf I324_inv Buffer
XI275 I331 I331_buf INV
XB275 I331_buf I331_inv Buffer
XI276 I332 I332_buf INV
XB276 I332_buf I332_inv Buffer
XI277 I333 I333_buf INV
XB277 I333_buf I333_inv Buffer
XI278 I334 I334_buf INV
XB278 I334_buf I334_inv Buffer
XI279 I341 I341_buf INV
XB279 I341_buf I341_inv Buffer
XI280 I342 I342_buf INV
XB280 I342_buf I342_inv Buffer
XI281 I343 I343_buf INV
XB281 I343_buf I343_inv Buffer
XI282 I344 I344_buf INV
XB282 I344_buf I344_inv Buffer
XI283 I351 I351_buf INV
XB283 I351_buf I351_inv Buffer
XI284 I352 I352_buf INV
XB284 I352_buf I352_inv Buffer
XI285 I353 I353_buf INV
XB285 I353_buf I353_inv Buffer
XI286 I354 I354_buf INV
XB286 I354_buf I354_inv Buffer
XI287 I361 I361_buf INV
XB287 I361_buf I361_inv Buffer
XI288 I362 I362_buf INV
XB288 I362_buf I362_inv Buffer
XI289 I363 I363_buf INV
XB289 I363_buf I363_inv Buffer
XI290 I364 I364_buf INV
XB290 I364_buf I364_inv Buffer
XI291 I371 I371_buf INV
XB291 I371_buf I371_inv Buffer
XI292 I372 I372_buf INV
XB292 I372_buf I372_inv Buffer
XI293 I373 I373_buf INV
XB293 I373_buf I373_inv Buffer
XI294 I374 I374_buf INV
XB294 I374_buf I374_inv Buffer
XI295 I381 I381_buf INV
XB295 I381_buf I381_inv Buffer
XI296 I382 I382_buf INV
XB296 I382_buf I382_inv Buffer
XI297 I383 I383_buf INV
XB297 I383_buf I383_inv Buffer
XI298 I384 I384_buf INV
XB298 I384_buf I384_inv Buffer
XI299 I391 I391_buf INV
XB299 I391_buf I391_inv Buffer
XI300 I392 I392_buf INV
XB300 I392_buf I392_inv Buffer
XI301 I393 I393_buf INV
XB301 I393_buf I393_inv Buffer
XI302 I394 I394_buf INV
XB302 I394_buf I394_inv Buffer
XI303 I3101 I3101_buf INV
XB303 I3101_buf I3101_inv Buffer
XI304 I3102 I3102_buf INV
XB304 I3102_buf I3102_inv Buffer
XI305 I3103 I3103_buf INV
XB305 I3103_buf I3103_inv Buffer
XI306 I3104 I3104_buf INV
XB306 I3104_buf I3104_inv Buffer
XI307 I3111 I3111_buf INV
XB307 I3111_buf I3111_inv Buffer
XI308 I3112 I3112_buf INV
XB308 I3112_buf I3112_inv Buffer
XI309 I3113 I3113_buf INV
XB309 I3113_buf I3113_inv Buffer
XI310 I3114 I3114_buf INV
XB310 I3114_buf I3114_inv Buffer
XI311 I3121 I3121_buf INV
XB311 I3121_buf I3121_inv Buffer
XI312 I3122 I3122_buf INV
XB312 I3122_buf I3122_inv Buffer
XI313 I3123 I3123_buf INV
XB313 I3123_buf I3123_inv Buffer
XI314 I3124 I3124_buf INV
XB314 I3124_buf I3124_inv Buffer
XI315 I3131 I3131_buf INV
XB315 I3131_buf I3131_inv Buffer
XI316 I3132 I3132_buf INV
XB316 I3132_buf I3132_inv Buffer
XI317 I3133 I3133_buf INV
XB317 I3133_buf I3133_inv Buffer
XI318 I3134 I3134_buf INV
XB318 I3134_buf I3134_inv Buffer
XI319 I3141 I3141_buf INV
XB319 I3141_buf I3141_inv Buffer
XI320 I3142 I3142_buf INV
XB320 I3142_buf I3142_inv Buffer
XI321 I3143 I3143_buf INV
XB321 I3143_buf I3143_inv Buffer
XI322 I3144 I3144_buf INV
XB322 I3144_buf I3144_inv Buffer
XI323 I3151 I3151_buf INV
XB323 I3151_buf I3151_inv Buffer
XI324 I3152 I3152_buf INV
XB324 I3152_buf I3152_inv Buffer
XI325 I3153 I3153_buf INV
XB325 I3153_buf I3153_inv Buffer
XI326 I3154 I3154_buf INV
XB326 I3154_buf I3154_inv Buffer
XI327 I3161 I3161_buf INV
XB327 I3161_buf I3161_inv Buffer
XI328 I3162 I3162_buf INV
XB328 I3162_buf I3162_inv Buffer
XI329 I3163 I3163_buf INV
XB329 I3163_buf I3163_inv Buffer
XI330 I3164 I3164_buf INV
XB330 I3164_buf I3164_inv Buffer
XI331 I3171 I3171_buf INV
XB331 I3171_buf I3171_inv Buffer
XI332 I3172 I3172_buf INV
XB332 I3172_buf I3172_inv Buffer
XI333 I3173 I3173_buf INV
XB333 I3173_buf I3173_inv Buffer
XI334 I3174 I3174_buf INV
XB334 I3174_buf I3174_inv Buffer
XI335 I3181 I3181_buf INV
XB335 I3181_buf I3181_inv Buffer
XI336 I3182 I3182_buf INV
XB336 I3182_buf I3182_inv Buffer
XI337 I3183 I3183_buf INV
XB337 I3183_buf I3183_inv Buffer
XI338 I3184 I3184_buf INV
XB338 I3184_buf I3184_inv Buffer
XI339 I3191 I3191_buf INV
XB339 I3191_buf I3191_inv Buffer
XI340 I3192 I3192_buf INV
XB340 I3192_buf I3192_inv Buffer
XI341 I3193 I3193_buf INV
XB341 I3193_buf I3193_inv Buffer
XI342 I3194 I3194_buf INV
XB342 I3194_buf I3194_inv Buffer
XI343 I3201 I3201_buf INV
XB343 I3201_buf I3201_inv Buffer
XI344 I3202 I3202_buf INV
XB344 I3202_buf I3202_inv Buffer
XI345 I3203 I3203_buf INV
XB345 I3203_buf I3203_inv Buffer
XI346 I3204 I3204_buf INV
XB346 I3204_buf I3204_inv Buffer
XI347 I3211 I3211_buf INV
XB347 I3211_buf I3211_inv Buffer
XI348 I3212 I3212_buf INV
XB348 I3212_buf I3212_inv Buffer
XI349 I3213 I3213_buf INV
XB349 I3213_buf I3213_inv Buffer
XI350 I3214 I3214_buf INV
XB350 I3214_buf I3214_inv Buffer
XI351 I3221 I3221_buf INV
XB351 I3221_buf I3221_inv Buffer
XI352 I3222 I3222_buf INV
XB352 I3222_buf I3222_inv Buffer
XI353 I3223 I3223_buf INV
XB353 I3223_buf I3223_inv Buffer
XI354 I3224 I3224_buf INV
XB354 I3224_buf I3224_inv Buffer
XI355 I3231 I3231_buf INV
XB355 I3231_buf I3231_inv Buffer
XI356 I3232 I3232_buf INV
XB356 I3232_buf I3232_inv Buffer
XI357 I3233 I3233_buf INV
XB357 I3233_buf I3233_inv Buffer
XI358 I3234 I3234_buf INV
XB358 I3234_buf I3234_inv Buffer
XI359 I3241 I3241_buf INV
XB359 I3241_buf I3241_inv Buffer
XI360 I3242 I3242_buf INV
XB360 I3242_buf I3242_inv Buffer
XI361 I3243 I3243_buf INV
XB361 I3243_buf I3243_inv Buffer
XI362 I3244 I3244_buf INV
XB362 I3244_buf I3244_inv Buffer
XI363 I3251 I3251_buf INV
XB363 I3251_buf I3251_inv Buffer
XI364 I3252 I3252_buf INV
XB364 I3252_buf I3252_inv Buffer
XI365 I3253 I3253_buf INV
XB365 I3253_buf I3253_inv Buffer
XI366 I3254 I3254_buf INV
XB366 I3254_buf I3254_inv Buffer
XI367 I3261 I3261_buf INV
XB367 I3261_buf I3261_inv Buffer
XI368 I3262 I3262_buf INV
XB368 I3262_buf I3262_inv Buffer
XI369 I3263 I3263_buf INV
XB369 I3263_buf I3263_inv Buffer
XI370 I3264 I3264_buf INV
XB370 I3264_buf I3264_inv Buffer
XI371 I3271 I3271_buf INV
XB371 I3271_buf I3271_inv Buffer
XI372 I3272 I3272_buf INV
XB372 I3272_buf I3272_inv Buffer
XI373 I3273 I3273_buf INV
XB373 I3273_buf I3273_inv Buffer
XI374 I3274 I3274_buf INV
XB374 I3274_buf I3274_inv Buffer
XI375 I3281 I3281_buf INV
XB375 I3281_buf I3281_inv Buffer
XI376 I3282 I3282_buf INV
XB376 I3282_buf I3282_inv Buffer
XI377 I3283 I3283_buf INV
XB377 I3283_buf I3283_inv Buffer
XI378 I3284 I3284_buf INV
XB378 I3284_buf I3284_inv Buffer
XI379 I3291 I3291_buf INV
XB379 I3291_buf I3291_inv Buffer
XI380 I3292 I3292_buf INV
XB380 I3292_buf I3292_inv Buffer
XI381 I3293 I3293_buf INV
XB381 I3293_buf I3293_inv Buffer
XI382 I3294 I3294_buf INV
XB382 I3294_buf I3294_inv Buffer
XI383 I3301 I3301_buf INV
XB383 I3301_buf I3301_inv Buffer
XI384 I3302 I3302_buf INV
XB384 I3302_buf I3302_inv Buffer
XI385 I3303 I3303_buf INV
XB385 I3303_buf I3303_inv Buffer
XI386 I3304 I3304_buf INV
XB386 I3304_buf I3304_inv Buffer
XI387 I3311 I3311_buf INV
XB387 I3311_buf I3311_inv Buffer
XI388 I3312 I3312_buf INV
XB388 I3312_buf I3312_inv Buffer
XI389 I3313 I3313_buf INV
XB389 I3313_buf I3313_inv Buffer
XI390 I3314 I3314_buf INV
XB390 I3314_buf I3314_inv Buffer
XI391 I3321 I3321_buf INV
XB391 I3321_buf I3321_inv Buffer
XI392 I3322 I3322_buf INV
XB392 I3322_buf I3322_inv Buffer
XI393 I3323 I3323_buf INV
XB393 I3323_buf I3323_inv Buffer
XI394 I3324 I3324_buf INV
XB394 I3324_buf I3324_inv Buffer
XI395 I411 I411_buf INV
XB395 I411_buf I411_inv Buffer
XI396 I412 I412_buf INV
XB396 I412_buf I412_inv Buffer
XI397 I413 I413_buf INV
XB397 I413_buf I413_inv Buffer
XI398 I414 I414_buf INV
XB398 I414_buf I414_inv Buffer
XI399 I421 I421_buf INV
XB399 I421_buf I421_inv Buffer
XI400 I422 I422_buf INV
XB400 I422_buf I422_inv Buffer
XI401 I423 I423_buf INV
XB401 I423_buf I423_inv Buffer
XI402 I424 I424_buf INV
XB402 I424_buf I424_inv Buffer
XI403 I431 I431_buf INV
XB403 I431_buf I431_inv Buffer
XI404 I432 I432_buf INV
XB404 I432_buf I432_inv Buffer
XI405 I433 I433_buf INV
XB405 I433_buf I433_inv Buffer
XI406 I434 I434_buf INV
XB406 I434_buf I434_inv Buffer
XI407 I441 I441_buf INV
XB407 I441_buf I441_inv Buffer
XI408 I442 I442_buf INV
XB408 I442_buf I442_inv Buffer
XI409 I443 I443_buf INV
XB409 I443_buf I443_inv Buffer
XI410 I444 I444_buf INV
XB410 I444_buf I444_inv Buffer
XI411 I451 I451_buf INV
XB411 I451_buf I451_inv Buffer
XI412 I452 I452_buf INV
XB412 I452_buf I452_inv Buffer
XI413 I453 I453_buf INV
XB413 I453_buf I453_inv Buffer
XI414 I454 I454_buf INV
XB414 I454_buf I454_inv Buffer
XI415 I461 I461_buf INV
XB415 I461_buf I461_inv Buffer
XI416 I462 I462_buf INV
XB416 I462_buf I462_inv Buffer
XI417 I463 I463_buf INV
XB417 I463_buf I463_inv Buffer
XI418 I464 I464_buf INV
XB418 I464_buf I464_inv Buffer
XI419 I471 I471_buf INV
XB419 I471_buf I471_inv Buffer
XI420 I472 I472_buf INV
XB420 I472_buf I472_inv Buffer
XI421 I473 I473_buf INV
XB421 I473_buf I473_inv Buffer
XI422 I474 I474_buf INV
XB422 I474_buf I474_inv Buffer
XI423 I481 I481_buf INV
XB423 I481_buf I481_inv Buffer
XI424 I482 I482_buf INV
XB424 I482_buf I482_inv Buffer
XI425 I483 I483_buf INV
XB425 I483_buf I483_inv Buffer
XI426 I484 I484_buf INV
XB426 I484_buf I484_inv Buffer
XI427 I491 I491_buf INV
XB427 I491_buf I491_inv Buffer
XI428 I492 I492_buf INV
XB428 I492_buf I492_inv Buffer
XI429 I493 I493_buf INV
XB429 I493_buf I493_inv Buffer
XI430 I494 I494_buf INV
XB430 I494_buf I494_inv Buffer
XI431 I4101 I4101_buf INV
XB431 I4101_buf I4101_inv Buffer
XI432 I4102 I4102_buf INV
XB432 I4102_buf I4102_inv Buffer
XI433 I4103 I4103_buf INV
XB433 I4103_buf I4103_inv Buffer
XI434 I4104 I4104_buf INV
XB434 I4104_buf I4104_inv Buffer
XI435 I4111 I4111_buf INV
XB435 I4111_buf I4111_inv Buffer
XI436 I4112 I4112_buf INV
XB436 I4112_buf I4112_inv Buffer
XI437 I4113 I4113_buf INV
XB437 I4113_buf I4113_inv Buffer
XI438 I4114 I4114_buf INV
XB438 I4114_buf I4114_inv Buffer
XI439 I4121 I4121_buf INV
XB439 I4121_buf I4121_inv Buffer
XI440 I4122 I4122_buf INV
XB440 I4122_buf I4122_inv Buffer
XI441 I4123 I4123_buf INV
XB441 I4123_buf I4123_inv Buffer
XI442 I4124 I4124_buf INV
XB442 I4124_buf I4124_inv Buffer
XI443 I4131 I4131_buf INV
XB443 I4131_buf I4131_inv Buffer
XI444 I4132 I4132_buf INV
XB444 I4132_buf I4132_inv Buffer
XI445 I4133 I4133_buf INV
XB445 I4133_buf I4133_inv Buffer
XI446 I4134 I4134_buf INV
XB446 I4134_buf I4134_inv Buffer
XI447 I4141 I4141_buf INV
XB447 I4141_buf I4141_inv Buffer
XI448 I4142 I4142_buf INV
XB448 I4142_buf I4142_inv Buffer
XI449 I4143 I4143_buf INV
XB449 I4143_buf I4143_inv Buffer
XI450 I4144 I4144_buf INV
XB450 I4144_buf I4144_inv Buffer
XI451 I4151 I4151_buf INV
XB451 I4151_buf I4151_inv Buffer
XI452 I4152 I4152_buf INV
XB452 I4152_buf I4152_inv Buffer
XI453 I4153 I4153_buf INV
XB453 I4153_buf I4153_inv Buffer
XI454 I4154 I4154_buf INV
XB454 I4154_buf I4154_inv Buffer
XI455 I4161 I4161_buf INV
XB455 I4161_buf I4161_inv Buffer
XI456 I4162 I4162_buf INV
XB456 I4162_buf I4162_inv Buffer
XI457 I4163 I4163_buf INV
XB457 I4163_buf I4163_inv Buffer
XI458 I4164 I4164_buf INV
XB458 I4164_buf I4164_inv Buffer
XI459 I4171 I4171_buf INV
XB459 I4171_buf I4171_inv Buffer
XI460 I4172 I4172_buf INV
XB460 I4172_buf I4172_inv Buffer
XI461 I4173 I4173_buf INV
XB461 I4173_buf I4173_inv Buffer
XI462 I4174 I4174_buf INV
XB462 I4174_buf I4174_inv Buffer
XI463 I4181 I4181_buf INV
XB463 I4181_buf I4181_inv Buffer
XI464 I4182 I4182_buf INV
XB464 I4182_buf I4182_inv Buffer
XI465 I4183 I4183_buf INV
XB465 I4183_buf I4183_inv Buffer
XI466 I4184 I4184_buf INV
XB466 I4184_buf I4184_inv Buffer
XI467 I4191 I4191_buf INV
XB467 I4191_buf I4191_inv Buffer
XI468 I4192 I4192_buf INV
XB468 I4192_buf I4192_inv Buffer
XI469 I4193 I4193_buf INV
XB469 I4193_buf I4193_inv Buffer
XI470 I4194 I4194_buf INV
XB470 I4194_buf I4194_inv Buffer
XI471 I4201 I4201_buf INV
XB471 I4201_buf I4201_inv Buffer
XI472 I4202 I4202_buf INV
XB472 I4202_buf I4202_inv Buffer
XI473 I4203 I4203_buf INV
XB473 I4203_buf I4203_inv Buffer
XI474 I4204 I4204_buf INV
XB474 I4204_buf I4204_inv Buffer
XI475 I4211 I4211_buf INV
XB475 I4211_buf I4211_inv Buffer
XI476 I4212 I4212_buf INV
XB476 I4212_buf I4212_inv Buffer
XI477 I4213 I4213_buf INV
XB477 I4213_buf I4213_inv Buffer
XI478 I4214 I4214_buf INV
XB478 I4214_buf I4214_inv Buffer
XI479 I4221 I4221_buf INV
XB479 I4221_buf I4221_inv Buffer
XI480 I4222 I4222_buf INV
XB480 I4222_buf I4222_inv Buffer
XI481 I4223 I4223_buf INV
XB481 I4223_buf I4223_inv Buffer
XI482 I4224 I4224_buf INV
XB482 I4224_buf I4224_inv Buffer
XI483 I4231 I4231_buf INV
XB483 I4231_buf I4231_inv Buffer
XI484 I4232 I4232_buf INV
XB484 I4232_buf I4232_inv Buffer
XI485 I4233 I4233_buf INV
XB485 I4233_buf I4233_inv Buffer
XI486 I4234 I4234_buf INV
XB486 I4234_buf I4234_inv Buffer
XI487 I4241 I4241_buf INV
XB487 I4241_buf I4241_inv Buffer
XI488 I4242 I4242_buf INV
XB488 I4242_buf I4242_inv Buffer
XI489 I4243 I4243_buf INV
XB489 I4243_buf I4243_inv Buffer
XI490 I4244 I4244_buf INV
XB490 I4244_buf I4244_inv Buffer
XI491 I4251 I4251_buf INV
XB491 I4251_buf I4251_inv Buffer
XI492 I4252 I4252_buf INV
XB492 I4252_buf I4252_inv Buffer
XI493 I4253 I4253_buf INV
XB493 I4253_buf I4253_inv Buffer
XI494 I4254 I4254_buf INV
XB494 I4254_buf I4254_inv Buffer
XI495 I4261 I4261_buf INV
XB495 I4261_buf I4261_inv Buffer
XI496 I4262 I4262_buf INV
XB496 I4262_buf I4262_inv Buffer
XI497 I4263 I4263_buf INV
XB497 I4263_buf I4263_inv Buffer
XI498 I4264 I4264_buf INV
XB498 I4264_buf I4264_inv Buffer
XI499 I4271 I4271_buf INV
XB499 I4271_buf I4271_inv Buffer
XI500 I4272 I4272_buf INV
XB500 I4272_buf I4272_inv Buffer
XI501 I4273 I4273_buf INV
XB501 I4273_buf I4273_inv Buffer
XI502 I4274 I4274_buf INV
XB502 I4274_buf I4274_inv Buffer
XI503 I4281 I4281_buf INV
XB503 I4281_buf I4281_inv Buffer
XI504 I4282 I4282_buf INV
XB504 I4282_buf I4282_inv Buffer
XI505 I4283 I4283_buf INV
XB505 I4283_buf I4283_inv Buffer
XI506 I4284 I4284_buf INV
XB506 I4284_buf I4284_inv Buffer
XI507 I4291 I4291_buf INV
XB507 I4291_buf I4291_inv Buffer
XI508 I4292 I4292_buf INV
XB508 I4292_buf I4292_inv Buffer
XI509 I4293 I4293_buf INV
XB509 I4293_buf I4293_inv Buffer
XI510 I4294 I4294_buf INV
XB510 I4294_buf I4294_inv Buffer
XI511 I4301 I4301_buf INV
XB511 I4301_buf I4301_inv Buffer
XI512 I4302 I4302_buf INV
XB512 I4302_buf I4302_inv Buffer
XI513 I4303 I4303_buf INV
XB513 I4303_buf I4303_inv Buffer
XI514 I4304 I4304_buf INV
XB514 I4304_buf I4304_inv Buffer
XI515 I4311 I4311_buf INV
XB515 I4311_buf I4311_inv Buffer
XI516 I4312 I4312_buf INV
XB516 I4312_buf I4312_inv Buffer
XI517 I4313 I4313_buf INV
XB517 I4313_buf I4313_inv Buffer
XI518 I4314 I4314_buf INV
XB518 I4314_buf I4314_inv Buffer
XI519 I4321 I4321_buf INV
XB519 I4321_buf I4321_inv Buffer
XI520 I4322 I4322_buf INV
XB520 I4322_buf I4322_inv Buffer
XI521 I4323 I4323_buf INV
XB521 I4323_buf I4323_inv Buffer
XI522 I4324 I4324_buf INV
XB522 I4324_buf I4324_inv Buffer



X1 I111_inv O_1_1_1 WL_1_1 BL BLB W_1_1_1 W_1_1_1_bar CIM_cell
X2 I112_inv O_1_1_2 WL_1_2 BL BLB W_1_1_2 W_1_1_2_bar CIM_cell
X3 I113_inv O_1_1_3 WL_1_3 BL BLB W_1_1_3 W_1_1_3_bar CIM_cell
X4 I114_inv O_1_1_4 WL_1_4 BL BLB W_1_1_4 W_1_1_4_bar CIM_cell
X5 I121_inv O_1_2_1 WL_1_1 BL BLB W_1_2_1 W_1_2_1_bar CIM_cell
X6 I122_inv O_1_2_2 WL_1_2 BL BLB W_1_2_2 W_1_2_2_bar CIM_cell
X7 I123_inv O_1_2_3 WL_1_3 BL BLB W_1_2_3 W_1_2_3_bar CIM_cell
X8 I124_inv O_1_2_4 WL_1_4 BL BLB W_1_2_4 W_1_2_4_bar CIM_cell
X9 I131_inv O_1_3_1 WL_1_1 BL BLB W_1_3_1 W_1_3_1_bar CIM_cell
X10 I132_inv O_1_3_2 WL_1_2 BL BLB W_1_3_2 W_1_3_2_bar CIM_cell
X11 I133_inv O_1_3_3 WL_1_3 BL BLB W_1_3_3 W_1_3_3_bar CIM_cell
X12 I134_inv O_1_3_4 WL_1_4 BL BLB W_1_3_4 W_1_3_4_bar CIM_cell
X13 I141_inv O_1_4_1 WL_1_1 BL BLB W_1_4_1 W_1_4_1_bar CIM_cell
X14 I142_inv O_1_4_2 WL_1_2 BL BLB W_1_4_2 W_1_4_2_bar CIM_cell
X15 I143_inv O_1_4_3 WL_1_3 BL BLB W_1_4_3 W_1_4_3_bar CIM_cell
X16 I144_inv O_1_4_4 WL_1_4 BL BLB W_1_4_4 W_1_4_4_bar CIM_cell
X17 I151_inv O_1_5_1 WL_1_1 BL BLB W_1_5_1 W_1_5_1_bar CIM_cell
X18 I152_inv O_1_5_2 WL_1_2 BL BLB W_1_5_2 W_1_5_2_bar CIM_cell
X19 I153_inv O_1_5_3 WL_1_3 BL BLB W_1_5_3 W_1_5_3_bar CIM_cell
X20 I154_inv O_1_5_4 WL_1_4 BL BLB W_1_5_4 W_1_5_4_bar CIM_cell
X21 I161_inv O_1_6_1 WL_1_1 BL BLB W_1_6_1 W_1_6_1_bar CIM_cell
X22 I162_inv O_1_6_2 WL_1_2 BL BLB W_1_6_2 W_1_6_2_bar CIM_cell
X23 I163_inv O_1_6_3 WL_1_3 BL BLB W_1_6_3 W_1_6_3_bar CIM_cell
X24 I164_inv O_1_6_4 WL_1_4 BL BLB W_1_6_4 W_1_6_4_bar CIM_cell
X25 I171_inv O_1_7_1 WL_1_1 BL BLB W_1_7_1 W_1_7_1_bar CIM_cell
X26 I172_inv O_1_7_2 WL_1_2 BL BLB W_1_7_2 W_1_7_2_bar CIM_cell
X27 I173_inv O_1_7_3 WL_1_3 BL BLB W_1_7_3 W_1_7_3_bar CIM_cell
X28 I174_inv O_1_7_4 WL_1_4 BL BLB W_1_7_4 W_1_7_4_bar CIM_cell
X29 I181_inv O_1_8_1 WL_1_1 BL BLB W_1_8_1 W_1_8_1_bar CIM_cell
X30 I182_inv O_1_8_2 WL_1_2 BL BLB W_1_8_2 W_1_8_2_bar CIM_cell
X31 I183_inv O_1_8_3 WL_1_3 BL BLB W_1_8_3 W_1_8_3_bar CIM_cell
X32 I184_inv O_1_8_4 WL_1_4 BL BLB W_1_8_4 W_1_8_4_bar CIM_cell
X33 I191_inv O_1_9_1 WL_1_1 BL BLB W_1_9_1 W_1_9_1_bar CIM_cell
X34 I192_inv O_1_9_2 WL_1_2 BL BLB W_1_9_2 W_1_9_2_bar CIM_cell
X35 I193_inv O_1_9_3 WL_1_3 BL BLB W_1_9_3 W_1_9_3_bar CIM_cell
X36 I194_inv O_1_9_4 WL_1_4 BL BLB W_1_9_4 W_1_9_4_bar CIM_cell
X37 I1101_inv O_1_10_1 WL_1_1 BL BLB W_1_10_1 W_1_10_1_bar CIM_cell
X38 I1102_inv O_1_10_2 WL_1_2 BL BLB W_1_10_2 W_1_10_2_bar CIM_cell
X39 I1103_inv O_1_10_3 WL_1_3 BL BLB W_1_10_3 W_1_10_3_bar CIM_cell
X40 I1104_inv O_1_10_4 WL_1_4 BL BLB W_1_10_4 W_1_10_4_bar CIM_cell
X41 I1111_inv O_1_11_1 WL_1_1 BL BLB W_1_11_1 W_1_11_1_bar CIM_cell
X42 I1112_inv O_1_11_2 WL_1_2 BL BLB W_1_11_2 W_1_11_2_bar CIM_cell
X43 I1113_inv O_1_11_3 WL_1_3 BL BLB W_1_11_3 W_1_11_3_bar CIM_cell
X44 I1114_inv O_1_11_4 WL_1_4 BL BLB W_1_11_4 W_1_11_4_bar CIM_cell
X45 I1121_inv O_1_12_1 WL_1_1 BL BLB W_1_12_1 W_1_12_1_bar CIM_cell
X46 I1122_inv O_1_12_2 WL_1_2 BL BLB W_1_12_2 W_1_12_2_bar CIM_cell
X47 I1123_inv O_1_12_3 WL_1_3 BL BLB W_1_12_3 W_1_12_3_bar CIM_cell
X48 I1124_inv O_1_12_4 WL_1_4 BL BLB W_1_12_4 W_1_12_4_bar CIM_cell
X49 I1131_inv O_1_13_1 WL_1_1 BL BLB W_1_13_1 W_1_13_1_bar CIM_cell
X50 I1132_inv O_1_13_2 WL_1_2 BL BLB W_1_13_2 W_1_13_2_bar CIM_cell
X51 I1133_inv O_1_13_3 WL_1_3 BL BLB W_1_13_3 W_1_13_3_bar CIM_cell
X52 I1134_inv O_1_13_4 WL_1_4 BL BLB W_1_13_4 W_1_13_4_bar CIM_cell
X53 I1141_inv O_1_14_1 WL_1_1 BL BLB W_1_14_1 W_1_14_1_bar CIM_cell
X54 I1142_inv O_1_14_2 WL_1_2 BL BLB W_1_14_2 W_1_14_2_bar CIM_cell
X55 I1143_inv O_1_14_3 WL_1_3 BL BLB W_1_14_3 W_1_14_3_bar CIM_cell
X56 I1144_inv O_1_14_4 WL_1_4 BL BLB W_1_14_4 W_1_14_4_bar CIM_cell
X57 I1151_inv O_1_15_1 WL_1_1 BL BLB W_1_15_1 W_1_15_1_bar CIM_cell
X58 I1152_inv O_1_15_2 WL_1_2 BL BLB W_1_15_2 W_1_15_2_bar CIM_cell
X59 I1153_inv O_1_15_3 WL_1_3 BL BLB W_1_15_3 W_1_15_3_bar CIM_cell
X60 I1154_inv O_1_15_4 WL_1_4 BL BLB W_1_15_4 W_1_15_4_bar CIM_cell
X61 I1161_inv O_1_16_1 WL_1_1 BL BLB W_1_16_1 W_1_16_1_bar CIM_cell
X62 I1162_inv O_1_16_2 WL_1_2 BL BLB W_1_16_2 W_1_16_2_bar CIM_cell
X63 I1163_inv O_1_16_3 WL_1_3 BL BLB W_1_16_3 W_1_16_3_bar CIM_cell
X64 I1164_inv O_1_16_4 WL_1_4 BL BLB W_1_16_4 W_1_16_4_bar CIM_cell
X65 I1171_inv O_1_17_1 WL_1_1 BL BLB W_1_17_1 W_1_17_1_bar CIM_cell
X66 I1172_inv O_1_17_2 WL_1_2 BL BLB W_1_17_2 W_1_17_2_bar CIM_cell
X67 I1173_inv O_1_17_3 WL_1_3 BL BLB W_1_17_3 W_1_17_3_bar CIM_cell
X68 I1174_inv O_1_17_4 WL_1_4 BL BLB W_1_17_4 W_1_17_4_bar CIM_cell
X69 I1181_inv O_1_18_1 WL_1_1 BL BLB W_1_18_1 W_1_18_1_bar CIM_cell
X70 I1182_inv O_1_18_2 WL_1_2 BL BLB W_1_18_2 W_1_18_2_bar CIM_cell
X71 I1183_inv O_1_18_3 WL_1_3 BL BLB W_1_18_3 W_1_18_3_bar CIM_cell
X72 I1184_inv O_1_18_4 WL_1_4 BL BLB W_1_18_4 W_1_18_4_bar CIM_cell
X73 I1191_inv O_1_19_1 WL_1_1 BL BLB W_1_19_1 W_1_19_1_bar CIM_cell
X74 I1192_inv O_1_19_2 WL_1_2 BL BLB W_1_19_2 W_1_19_2_bar CIM_cell
X75 I1193_inv O_1_19_3 WL_1_3 BL BLB W_1_19_3 W_1_19_3_bar CIM_cell
X76 I1194_inv O_1_19_4 WL_1_4 BL BLB W_1_19_4 W_1_19_4_bar CIM_cell
X77 I1201_inv O_1_20_1 WL_1_1 BL BLB W_1_20_1 W_1_20_1_bar CIM_cell
X78 I1202_inv O_1_20_2 WL_1_2 BL BLB W_1_20_2 W_1_20_2_bar CIM_cell
X79 I1203_inv O_1_20_3 WL_1_3 BL BLB W_1_20_3 W_1_20_3_bar CIM_cell
X80 I1204_inv O_1_20_4 WL_1_4 BL BLB W_1_20_4 W_1_20_4_bar CIM_cell
X81 I1211_inv O_1_21_1 WL_1_1 BL BLB W_1_21_1 W_1_21_1_bar CIM_cell
X82 I1212_inv O_1_21_2 WL_1_2 BL BLB W_1_21_2 W_1_21_2_bar CIM_cell
X83 I1213_inv O_1_21_3 WL_1_3 BL BLB W_1_21_3 W_1_21_3_bar CIM_cell
X84 I1214_inv O_1_21_4 WL_1_4 BL BLB W_1_21_4 W_1_21_4_bar CIM_cell
X85 I1221_inv O_1_22_1 WL_1_1 BL BLB W_1_22_1 W_1_22_1_bar CIM_cell
X86 I1222_inv O_1_22_2 WL_1_2 BL BLB W_1_22_2 W_1_22_2_bar CIM_cell
X87 I1223_inv O_1_22_3 WL_1_3 BL BLB W_1_22_3 W_1_22_3_bar CIM_cell
X88 I1224_inv O_1_22_4 WL_1_4 BL BLB W_1_22_4 W_1_22_4_bar CIM_cell
X89 I1231_inv O_1_23_1 WL_1_1 BL BLB W_1_23_1 W_1_23_1_bar CIM_cell
X90 I1232_inv O_1_23_2 WL_1_2 BL BLB W_1_23_2 W_1_23_2_bar CIM_cell
X91 I1233_inv O_1_23_3 WL_1_3 BL BLB W_1_23_3 W_1_23_3_bar CIM_cell
X92 I1234_inv O_1_23_4 WL_1_4 BL BLB W_1_23_4 W_1_23_4_bar CIM_cell
X93 I1241_inv O_1_24_1 WL_1_1 BL BLB W_1_24_1 W_1_24_1_bar CIM_cell
X94 I1242_inv O_1_24_2 WL_1_2 BL BLB W_1_24_2 W_1_24_2_bar CIM_cell
X95 I1243_inv O_1_24_3 WL_1_3 BL BLB W_1_24_3 W_1_24_3_bar CIM_cell
X96 I1244_inv O_1_24_4 WL_1_4 BL BLB W_1_24_4 W_1_24_4_bar CIM_cell
X97 I1251_inv O_1_25_1 WL_1_1 BL BLB W_1_25_1 W_1_25_1_bar CIM_cell
X98 I1252_inv O_1_25_2 WL_1_2 BL BLB W_1_25_2 W_1_25_2_bar CIM_cell
X99 I1253_inv O_1_25_3 WL_1_3 BL BLB W_1_25_3 W_1_25_3_bar CIM_cell
X100 I1254_inv O_1_25_4 WL_1_4 BL BLB W_1_25_4 W_1_25_4_bar CIM_cell
X101 I1261_inv O_1_26_1 WL_1_1 BL BLB W_1_26_1 W_1_26_1_bar CIM_cell
X102 I1262_inv O_1_26_2 WL_1_2 BL BLB W_1_26_2 W_1_26_2_bar CIM_cell
X103 I1263_inv O_1_26_3 WL_1_3 BL BLB W_1_26_3 W_1_26_3_bar CIM_cell
X104 I1264_inv O_1_26_4 WL_1_4 BL BLB W_1_26_4 W_1_26_4_bar CIM_cell
X105 I1271_inv O_1_27_1 WL_1_1 BL BLB W_1_27_1 W_1_27_1_bar CIM_cell
X106 I1272_inv O_1_27_2 WL_1_2 BL BLB W_1_27_2 W_1_27_2_bar CIM_cell
X107 I1273_inv O_1_27_3 WL_1_3 BL BLB W_1_27_3 W_1_27_3_bar CIM_cell
X108 I1274_inv O_1_27_4 WL_1_4 BL BLB W_1_27_4 W_1_27_4_bar CIM_cell
X109 I1281_inv O_1_28_1 WL_1_1 BL BLB W_1_28_1 W_1_28_1_bar CIM_cell
X110 I1282_inv O_1_28_2 WL_1_2 BL BLB W_1_28_2 W_1_28_2_bar CIM_cell
X111 I1283_inv O_1_28_3 WL_1_3 BL BLB W_1_28_3 W_1_28_3_bar CIM_cell
X112 I1284_inv O_1_28_4 WL_1_4 BL BLB W_1_28_4 W_1_28_4_bar CIM_cell
X113 I1291_inv O_1_29_1 WL_1_1 BL BLB W_1_29_1 W_1_29_1_bar CIM_cell
X114 I1292_inv O_1_29_2 WL_1_2 BL BLB W_1_29_2 W_1_29_2_bar CIM_cell
X115 I1293_inv O_1_29_3 WL_1_3 BL BLB W_1_29_3 W_1_29_3_bar CIM_cell
X116 I1294_inv O_1_29_4 WL_1_4 BL BLB W_1_29_4 W_1_29_4_bar CIM_cell
X117 I1301_inv O_1_30_1 WL_1_1 BL BLB W_1_30_1 W_1_30_1_bar CIM_cell
X118 I1302_inv O_1_30_2 WL_1_2 BL BLB W_1_30_2 W_1_30_2_bar CIM_cell
X119 I1303_inv O_1_30_3 WL_1_3 BL BLB W_1_30_3 W_1_30_3_bar CIM_cell
X120 I1304_inv O_1_30_4 WL_1_4 BL BLB W_1_30_4 W_1_30_4_bar CIM_cell
X121 I1311_inv O_1_31_1 WL_1_1 BL BLB W_1_31_1 W_1_31_1_bar CIM_cell
X122 I1312_inv O_1_31_2 WL_1_2 BL BLB W_1_31_2 W_1_31_2_bar CIM_cell
X123 I1313_inv O_1_31_3 WL_1_3 BL BLB W_1_31_3 W_1_31_3_bar CIM_cell
X124 I1314_inv O_1_31_4 WL_1_4 BL BLB W_1_31_4 W_1_31_4_bar CIM_cell
X125 I1321_inv O_1_32_1 WL_1_1 BL BLB W_1_32_1 W_1_32_1_bar CIM_cell
X126 I1322_inv O_1_32_2 WL_1_2 BL BLB W_1_32_2 W_1_32_2_bar CIM_cell
X127 I1323_inv O_1_32_3 WL_1_3 BL BLB W_1_32_3 W_1_32_3_bar CIM_cell
X128 I1324_inv O_1_32_4 WL_1_4 BL BLB W_1_32_4 W_1_32_4_bar CIM_cell
X129 I211_inv O_2_1_1 WL_2_1 BL BLB W_2_1_1 W_2_1_1_bar CIM_cell
X130 I212_inv O_2_1_2 WL_2_2 BL BLB W_2_1_2 W_2_1_2_bar CIM_cell
X131 I213_inv O_2_1_3 WL_2_3 BL BLB W_2_1_3 W_2_1_3_bar CIM_cell
X132 I214_inv O_2_1_4 WL_2_4 BL BLB W_2_1_4 W_2_1_4_bar CIM_cell
X133 I221_inv O_2_2_1 WL_2_1 BL BLB W_2_2_1 W_2_2_1_bar CIM_cell
X134 I222_inv O_2_2_2 WL_2_2 BL BLB W_2_2_2 W_2_2_2_bar CIM_cell
X135 I223_inv O_2_2_3 WL_2_3 BL BLB W_2_2_3 W_2_2_3_bar CIM_cell
X136 I224_inv O_2_2_4 WL_2_4 BL BLB W_2_2_4 W_2_2_4_bar CIM_cell
X137 I231_inv O_2_3_1 WL_2_1 BL BLB W_2_3_1 W_2_3_1_bar CIM_cell
X138 I232_inv O_2_3_2 WL_2_2 BL BLB W_2_3_2 W_2_3_2_bar CIM_cell
X139 I233_inv O_2_3_3 WL_2_3 BL BLB W_2_3_3 W_2_3_3_bar CIM_cell
X140 I234_inv O_2_3_4 WL_2_4 BL BLB W_2_3_4 W_2_3_4_bar CIM_cell
X141 I241_inv O_2_4_1 WL_2_1 BL BLB W_2_4_1 W_2_4_1_bar CIM_cell
X142 I242_inv O_2_4_2 WL_2_2 BL BLB W_2_4_2 W_2_4_2_bar CIM_cell
X143 I243_inv O_2_4_3 WL_2_3 BL BLB W_2_4_3 W_2_4_3_bar CIM_cell
X144 I244_inv O_2_4_4 WL_2_4 BL BLB W_2_4_4 W_2_4_4_bar CIM_cell
X145 I251_inv O_2_5_1 WL_2_1 BL BLB W_2_5_1 W_2_5_1_bar CIM_cell
X146 I252_inv O_2_5_2 WL_2_2 BL BLB W_2_5_2 W_2_5_2_bar CIM_cell
X147 I253_inv O_2_5_3 WL_2_3 BL BLB W_2_5_3 W_2_5_3_bar CIM_cell
X148 I254_inv O_2_5_4 WL_2_4 BL BLB W_2_5_4 W_2_5_4_bar CIM_cell
X149 I261_inv O_2_6_1 WL_2_1 BL BLB W_2_6_1 W_2_6_1_bar CIM_cell
X150 I262_inv O_2_6_2 WL_2_2 BL BLB W_2_6_2 W_2_6_2_bar CIM_cell
X151 I263_inv O_2_6_3 WL_2_3 BL BLB W_2_6_3 W_2_6_3_bar CIM_cell
X152 I264_inv O_2_6_4 WL_2_4 BL BLB W_2_6_4 W_2_6_4_bar CIM_cell
X153 I271_inv O_2_7_1 WL_2_1 BL BLB W_2_7_1 W_2_7_1_bar CIM_cell
X154 I272_inv O_2_7_2 WL_2_2 BL BLB W_2_7_2 W_2_7_2_bar CIM_cell
X155 I273_inv O_2_7_3 WL_2_3 BL BLB W_2_7_3 W_2_7_3_bar CIM_cell
X156 I274_inv O_2_7_4 WL_2_4 BL BLB W_2_7_4 W_2_7_4_bar CIM_cell
X157 I281_inv O_2_8_1 WL_2_1 BL BLB W_2_8_1 W_2_8_1_bar CIM_cell
X158 I282_inv O_2_8_2 WL_2_2 BL BLB W_2_8_2 W_2_8_2_bar CIM_cell
X159 I283_inv O_2_8_3 WL_2_3 BL BLB W_2_8_3 W_2_8_3_bar CIM_cell
X160 I284_inv O_2_8_4 WL_2_4 BL BLB W_2_8_4 W_2_8_4_bar CIM_cell
X161 I291_inv O_2_9_1 WL_2_1 BL BLB W_2_9_1 W_2_9_1_bar CIM_cell
X162 I292_inv O_2_9_2 WL_2_2 BL BLB W_2_9_2 W_2_9_2_bar CIM_cell
X163 I293_inv O_2_9_3 WL_2_3 BL BLB W_2_9_3 W_2_9_3_bar CIM_cell
X164 I294_inv O_2_9_4 WL_2_4 BL BLB W_2_9_4 W_2_9_4_bar CIM_cell
X165 I2101_inv O_2_10_1 WL_2_1 BL BLB W_2_10_1 W_2_10_1_bar CIM_cell
X166 I2102_inv O_2_10_2 WL_2_2 BL BLB W_2_10_2 W_2_10_2_bar CIM_cell
X167 I2103_inv O_2_10_3 WL_2_3 BL BLB W_2_10_3 W_2_10_3_bar CIM_cell
X168 I2104_inv O_2_10_4 WL_2_4 BL BLB W_2_10_4 W_2_10_4_bar CIM_cell
X169 I2111_inv O_2_11_1 WL_2_1 BL BLB W_2_11_1 W_2_11_1_bar CIM_cell
X170 I2112_inv O_2_11_2 WL_2_2 BL BLB W_2_11_2 W_2_11_2_bar CIM_cell
X171 I2113_inv O_2_11_3 WL_2_3 BL BLB W_2_11_3 W_2_11_3_bar CIM_cell
X172 I2114_inv O_2_11_4 WL_2_4 BL BLB W_2_11_4 W_2_11_4_bar CIM_cell
X173 I2121_inv O_2_12_1 WL_2_1 BL BLB W_2_12_1 W_2_12_1_bar CIM_cell
X174 I2122_inv O_2_12_2 WL_2_2 BL BLB W_2_12_2 W_2_12_2_bar CIM_cell
X175 I2123_inv O_2_12_3 WL_2_3 BL BLB W_2_12_3 W_2_12_3_bar CIM_cell
X176 I2124_inv O_2_12_4 WL_2_4 BL BLB W_2_12_4 W_2_12_4_bar CIM_cell
X177 I2131_inv O_2_13_1 WL_2_1 BL BLB W_2_13_1 W_2_13_1_bar CIM_cell
X178 I2132_inv O_2_13_2 WL_2_2 BL BLB W_2_13_2 W_2_13_2_bar CIM_cell
X179 I2133_inv O_2_13_3 WL_2_3 BL BLB W_2_13_3 W_2_13_3_bar CIM_cell
X180 I2134_inv O_2_13_4 WL_2_4 BL BLB W_2_13_4 W_2_13_4_bar CIM_cell
X181 I2141_inv O_2_14_1 WL_2_1 BL BLB W_2_14_1 W_2_14_1_bar CIM_cell
X182 I2142_inv O_2_14_2 WL_2_2 BL BLB W_2_14_2 W_2_14_2_bar CIM_cell
X183 I2143_inv O_2_14_3 WL_2_3 BL BLB W_2_14_3 W_2_14_3_bar CIM_cell
X184 I2144_inv O_2_14_4 WL_2_4 BL BLB W_2_14_4 W_2_14_4_bar CIM_cell
X185 I2151_inv O_2_15_1 WL_2_1 BL BLB W_2_15_1 W_2_15_1_bar CIM_cell
X186 I2152_inv O_2_15_2 WL_2_2 BL BLB W_2_15_2 W_2_15_2_bar CIM_cell
X187 I2153_inv O_2_15_3 WL_2_3 BL BLB W_2_15_3 W_2_15_3_bar CIM_cell
X188 I2154_inv O_2_15_4 WL_2_4 BL BLB W_2_15_4 W_2_15_4_bar CIM_cell
X189 I2161_inv O_2_16_1 WL_2_1 BL BLB W_2_16_1 W_2_16_1_bar CIM_cell
X190 I2162_inv O_2_16_2 WL_2_2 BL BLB W_2_16_2 W_2_16_2_bar CIM_cell
X191 I2163_inv O_2_16_3 WL_2_3 BL BLB W_2_16_3 W_2_16_3_bar CIM_cell
X192 I2164_inv O_2_16_4 WL_2_4 BL BLB W_2_16_4 W_2_16_4_bar CIM_cell
X193 I2171_inv O_2_17_1 WL_2_1 BL BLB W_2_17_1 W_2_17_1_bar CIM_cell
X194 I2172_inv O_2_17_2 WL_2_2 BL BLB W_2_17_2 W_2_17_2_bar CIM_cell
X195 I2173_inv O_2_17_3 WL_2_3 BL BLB W_2_17_3 W_2_17_3_bar CIM_cell
X196 I2174_inv O_2_17_4 WL_2_4 BL BLB W_2_17_4 W_2_17_4_bar CIM_cell
X197 I2181_inv O_2_18_1 WL_2_1 BL BLB W_2_18_1 W_2_18_1_bar CIM_cell
X198 I2182_inv O_2_18_2 WL_2_2 BL BLB W_2_18_2 W_2_18_2_bar CIM_cell
X199 I2183_inv O_2_18_3 WL_2_3 BL BLB W_2_18_3 W_2_18_3_bar CIM_cell
X200 I2184_inv O_2_18_4 WL_2_4 BL BLB W_2_18_4 W_2_18_4_bar CIM_cell
X201 I2191_inv O_2_19_1 WL_2_1 BL BLB W_2_19_1 W_2_19_1_bar CIM_cell
X202 I2192_inv O_2_19_2 WL_2_2 BL BLB W_2_19_2 W_2_19_2_bar CIM_cell
X203 I2193_inv O_2_19_3 WL_2_3 BL BLB W_2_19_3 W_2_19_3_bar CIM_cell
X204 I2194_inv O_2_19_4 WL_2_4 BL BLB W_2_19_4 W_2_19_4_bar CIM_cell
X205 I2201_inv O_2_20_1 WL_2_1 BL BLB W_2_20_1 W_2_20_1_bar CIM_cell
X206 I2202_inv O_2_20_2 WL_2_2 BL BLB W_2_20_2 W_2_20_2_bar CIM_cell
X207 I2203_inv O_2_20_3 WL_2_3 BL BLB W_2_20_3 W_2_20_3_bar CIM_cell
X208 I2204_inv O_2_20_4 WL_2_4 BL BLB W_2_20_4 W_2_20_4_bar CIM_cell
X209 I2211_inv O_2_21_1 WL_2_1 BL BLB W_2_21_1 W_2_21_1_bar CIM_cell
X210 I2212_inv O_2_21_2 WL_2_2 BL BLB W_2_21_2 W_2_21_2_bar CIM_cell
X211 I2213_inv O_2_21_3 WL_2_3 BL BLB W_2_21_3 W_2_21_3_bar CIM_cell
X212 I2214_inv O_2_21_4 WL_2_4 BL BLB W_2_21_4 W_2_21_4_bar CIM_cell
X213 I2221_inv O_2_22_1 WL_2_1 BL BLB W_2_22_1 W_2_22_1_bar CIM_cell
X214 I2222_inv O_2_22_2 WL_2_2 BL BLB W_2_22_2 W_2_22_2_bar CIM_cell
X215 I2223_inv O_2_22_3 WL_2_3 BL BLB W_2_22_3 W_2_22_3_bar CIM_cell
X216 I2224_inv O_2_22_4 WL_2_4 BL BLB W_2_22_4 W_2_22_4_bar CIM_cell
X217 I2231_inv O_2_23_1 WL_2_1 BL BLB W_2_23_1 W_2_23_1_bar CIM_cell
X218 I2232_inv O_2_23_2 WL_2_2 BL BLB W_2_23_2 W_2_23_2_bar CIM_cell
X219 I2233_inv O_2_23_3 WL_2_3 BL BLB W_2_23_3 W_2_23_3_bar CIM_cell
X220 I2234_inv O_2_23_4 WL_2_4 BL BLB W_2_23_4 W_2_23_4_bar CIM_cell
X221 I2241_inv O_2_24_1 WL_2_1 BL BLB W_2_24_1 W_2_24_1_bar CIM_cell
X222 I2242_inv O_2_24_2 WL_2_2 BL BLB W_2_24_2 W_2_24_2_bar CIM_cell
X223 I2243_inv O_2_24_3 WL_2_3 BL BLB W_2_24_3 W_2_24_3_bar CIM_cell
X224 I2244_inv O_2_24_4 WL_2_4 BL BLB W_2_24_4 W_2_24_4_bar CIM_cell
X225 I2251_inv O_2_25_1 WL_2_1 BL BLB W_2_25_1 W_2_25_1_bar CIM_cell
X226 I2252_inv O_2_25_2 WL_2_2 BL BLB W_2_25_2 W_2_25_2_bar CIM_cell
X227 I2253_inv O_2_25_3 WL_2_3 BL BLB W_2_25_3 W_2_25_3_bar CIM_cell
X228 I2254_inv O_2_25_4 WL_2_4 BL BLB W_2_25_4 W_2_25_4_bar CIM_cell
X229 I2261_inv O_2_26_1 WL_2_1 BL BLB W_2_26_1 W_2_26_1_bar CIM_cell
X230 I2262_inv O_2_26_2 WL_2_2 BL BLB W_2_26_2 W_2_26_2_bar CIM_cell
X231 I2263_inv O_2_26_3 WL_2_3 BL BLB W_2_26_3 W_2_26_3_bar CIM_cell
X232 I2264_inv O_2_26_4 WL_2_4 BL BLB W_2_26_4 W_2_26_4_bar CIM_cell
X233 I2271_inv O_2_27_1 WL_2_1 BL BLB W_2_27_1 W_2_27_1_bar CIM_cell
X234 I2272_inv O_2_27_2 WL_2_2 BL BLB W_2_27_2 W_2_27_2_bar CIM_cell
X235 I2273_inv O_2_27_3 WL_2_3 BL BLB W_2_27_3 W_2_27_3_bar CIM_cell
X236 I2274_inv O_2_27_4 WL_2_4 BL BLB W_2_27_4 W_2_27_4_bar CIM_cell
X237 I2281_inv O_2_28_1 WL_2_1 BL BLB W_2_28_1 W_2_28_1_bar CIM_cell
X238 I2282_inv O_2_28_2 WL_2_2 BL BLB W_2_28_2 W_2_28_2_bar CIM_cell
X239 I2283_inv O_2_28_3 WL_2_3 BL BLB W_2_28_3 W_2_28_3_bar CIM_cell
X240 I2284_inv O_2_28_4 WL_2_4 BL BLB W_2_28_4 W_2_28_4_bar CIM_cell
X241 I2291_inv O_2_29_1 WL_2_1 BL BLB W_2_29_1 W_2_29_1_bar CIM_cell
X242 I2292_inv O_2_29_2 WL_2_2 BL BLB W_2_29_2 W_2_29_2_bar CIM_cell
X243 I2293_inv O_2_29_3 WL_2_3 BL BLB W_2_29_3 W_2_29_3_bar CIM_cell
X244 I2294_inv O_2_29_4 WL_2_4 BL BLB W_2_29_4 W_2_29_4_bar CIM_cell
X245 I2301_inv O_2_30_1 WL_2_1 BL BLB W_2_30_1 W_2_30_1_bar CIM_cell
X246 I2302_inv O_2_30_2 WL_2_2 BL BLB W_2_30_2 W_2_30_2_bar CIM_cell
X247 I2303_inv O_2_30_3 WL_2_3 BL BLB W_2_30_3 W_2_30_3_bar CIM_cell
X248 I2304_inv O_2_30_4 WL_2_4 BL BLB W_2_30_4 W_2_30_4_bar CIM_cell
X249 I2311_inv O_2_31_1 WL_2_1 BL BLB W_2_31_1 W_2_31_1_bar CIM_cell
X250 I2312_inv O_2_31_2 WL_2_2 BL BLB W_2_31_2 W_2_31_2_bar CIM_cell
X251 I2313_inv O_2_31_3 WL_2_3 BL BLB W_2_31_3 W_2_31_3_bar CIM_cell
X252 I2314_inv O_2_31_4 WL_2_4 BL BLB W_2_31_4 W_2_31_4_bar CIM_cell
X253 I2321_inv O_2_32_1 WL_2_1 BL BLB W_2_32_1 W_2_32_1_bar CIM_cell
X254 I2322_inv O_2_32_2 WL_2_2 BL BLB W_2_32_2 W_2_32_2_bar CIM_cell
X255 I2323_inv O_2_32_3 WL_2_3 BL BLB W_2_32_3 W_2_32_3_bar CIM_cell
X256 I2324_inv O_2_32_4 WL_2_4 BL BLB W_2_32_4 W_2_32_4_bar CIM_cell
X257 I311_inv O_3_1_1 WL_3_1 BL BLB W_3_1_1 W_3_1_1_bar CIM_cell
X258 I312_inv O_3_1_2 WL_3_2 BL BLB W_3_1_2 W_3_1_2_bar CIM_cell
X259 I313_inv O_3_1_3 WL_3_3 BL BLB W_3_1_3 W_3_1_3_bar CIM_cell
X260 I314_inv O_3_1_4 WL_3_4 BL BLB W_3_1_4 W_3_1_4_bar CIM_cell
X261 I321_inv O_3_2_1 WL_3_1 BL BLB W_3_2_1 W_3_2_1_bar CIM_cell
X262 I322_inv O_3_2_2 WL_3_2 BL BLB W_3_2_2 W_3_2_2_bar CIM_cell
X263 I323_inv O_3_2_3 WL_3_3 BL BLB W_3_2_3 W_3_2_3_bar CIM_cell
X264 I324_inv O_3_2_4 WL_3_4 BL BLB W_3_2_4 W_3_2_4_bar CIM_cell
X265 I331_inv O_3_3_1 WL_3_1 BL BLB W_3_3_1 W_3_3_1_bar CIM_cell
X266 I332_inv O_3_3_2 WL_3_2 BL BLB W_3_3_2 W_3_3_2_bar CIM_cell
X267 I333_inv O_3_3_3 WL_3_3 BL BLB W_3_3_3 W_3_3_3_bar CIM_cell
X268 I334_inv O_3_3_4 WL_3_4 BL BLB W_3_3_4 W_3_3_4_bar CIM_cell
X269 I341_inv O_3_4_1 WL_3_1 BL BLB W_3_4_1 W_3_4_1_bar CIM_cell
X270 I342_inv O_3_4_2 WL_3_2 BL BLB W_3_4_2 W_3_4_2_bar CIM_cell
X271 I343_inv O_3_4_3 WL_3_3 BL BLB W_3_4_3 W_3_4_3_bar CIM_cell
X272 I344_inv O_3_4_4 WL_3_4 BL BLB W_3_4_4 W_3_4_4_bar CIM_cell
X273 I351_inv O_3_5_1 WL_3_1 BL BLB W_3_5_1 W_3_5_1_bar CIM_cell
X274 I352_inv O_3_5_2 WL_3_2 BL BLB W_3_5_2 W_3_5_2_bar CIM_cell
X275 I353_inv O_3_5_3 WL_3_3 BL BLB W_3_5_3 W_3_5_3_bar CIM_cell
X276 I354_inv O_3_5_4 WL_3_4 BL BLB W_3_5_4 W_3_5_4_bar CIM_cell
X277 I361_inv O_3_6_1 WL_3_1 BL BLB W_3_6_1 W_3_6_1_bar CIM_cell
X278 I362_inv O_3_6_2 WL_3_2 BL BLB W_3_6_2 W_3_6_2_bar CIM_cell
X279 I363_inv O_3_6_3 WL_3_3 BL BLB W_3_6_3 W_3_6_3_bar CIM_cell
X280 I364_inv O_3_6_4 WL_3_4 BL BLB W_3_6_4 W_3_6_4_bar CIM_cell
X281 I371_inv O_3_7_1 WL_3_1 BL BLB W_3_7_1 W_3_7_1_bar CIM_cell
X282 I372_inv O_3_7_2 WL_3_2 BL BLB W_3_7_2 W_3_7_2_bar CIM_cell
X283 I373_inv O_3_7_3 WL_3_3 BL BLB W_3_7_3 W_3_7_3_bar CIM_cell
X284 I374_inv O_3_7_4 WL_3_4 BL BLB W_3_7_4 W_3_7_4_bar CIM_cell
X285 I381_inv O_3_8_1 WL_3_1 BL BLB W_3_8_1 W_3_8_1_bar CIM_cell
X286 I382_inv O_3_8_2 WL_3_2 BL BLB W_3_8_2 W_3_8_2_bar CIM_cell
X287 I383_inv O_3_8_3 WL_3_3 BL BLB W_3_8_3 W_3_8_3_bar CIM_cell
X288 I384_inv O_3_8_4 WL_3_4 BL BLB W_3_8_4 W_3_8_4_bar CIM_cell
X289 I391_inv O_3_9_1 WL_3_1 BL BLB W_3_9_1 W_3_9_1_bar CIM_cell
X290 I392_inv O_3_9_2 WL_3_2 BL BLB W_3_9_2 W_3_9_2_bar CIM_cell
X291 I393_inv O_3_9_3 WL_3_3 BL BLB W_3_9_3 W_3_9_3_bar CIM_cell
X292 I394_inv O_3_9_4 WL_3_4 BL BLB W_3_9_4 W_3_9_4_bar CIM_cell
X293 I3101_inv O_3_10_1 WL_3_1 BL BLB W_3_10_1 W_3_10_1_bar CIM_cell
X294 I3102_inv O_3_10_2 WL_3_2 BL BLB W_3_10_2 W_3_10_2_bar CIM_cell
X295 I3103_inv O_3_10_3 WL_3_3 BL BLB W_3_10_3 W_3_10_3_bar CIM_cell
X296 I3104_inv O_3_10_4 WL_3_4 BL BLB W_3_10_4 W_3_10_4_bar CIM_cell
X297 I3111_inv O_3_11_1 WL_3_1 BL BLB W_3_11_1 W_3_11_1_bar CIM_cell
X298 I3112_inv O_3_11_2 WL_3_2 BL BLB W_3_11_2 W_3_11_2_bar CIM_cell
X299 I3113_inv O_3_11_3 WL_3_3 BL BLB W_3_11_3 W_3_11_3_bar CIM_cell
X300 I3114_inv O_3_11_4 WL_3_4 BL BLB W_3_11_4 W_3_11_4_bar CIM_cell
X301 I3121_inv O_3_12_1 WL_3_1 BL BLB W_3_12_1 W_3_12_1_bar CIM_cell
X302 I3122_inv O_3_12_2 WL_3_2 BL BLB W_3_12_2 W_3_12_2_bar CIM_cell
X303 I3123_inv O_3_12_3 WL_3_3 BL BLB W_3_12_3 W_3_12_3_bar CIM_cell
X304 I3124_inv O_3_12_4 WL_3_4 BL BLB W_3_12_4 W_3_12_4_bar CIM_cell
X305 I3131_inv O_3_13_1 WL_3_1 BL BLB W_3_13_1 W_3_13_1_bar CIM_cell
X306 I3132_inv O_3_13_2 WL_3_2 BL BLB W_3_13_2 W_3_13_2_bar CIM_cell
X307 I3133_inv O_3_13_3 WL_3_3 BL BLB W_3_13_3 W_3_13_3_bar CIM_cell
X308 I3134_inv O_3_13_4 WL_3_4 BL BLB W_3_13_4 W_3_13_4_bar CIM_cell
X309 I3141_inv O_3_14_1 WL_3_1 BL BLB W_3_14_1 W_3_14_1_bar CIM_cell
X310 I3142_inv O_3_14_2 WL_3_2 BL BLB W_3_14_2 W_3_14_2_bar CIM_cell
X311 I3143_inv O_3_14_3 WL_3_3 BL BLB W_3_14_3 W_3_14_3_bar CIM_cell
X312 I3144_inv O_3_14_4 WL_3_4 BL BLB W_3_14_4 W_3_14_4_bar CIM_cell
X313 I3151_inv O_3_15_1 WL_3_1 BL BLB W_3_15_1 W_3_15_1_bar CIM_cell
X314 I3152_inv O_3_15_2 WL_3_2 BL BLB W_3_15_2 W_3_15_2_bar CIM_cell
X315 I3153_inv O_3_15_3 WL_3_3 BL BLB W_3_15_3 W_3_15_3_bar CIM_cell
X316 I3154_inv O_3_15_4 WL_3_4 BL BLB W_3_15_4 W_3_15_4_bar CIM_cell
X317 I3161_inv O_3_16_1 WL_3_1 BL BLB W_3_16_1 W_3_16_1_bar CIM_cell
X318 I3162_inv O_3_16_2 WL_3_2 BL BLB W_3_16_2 W_3_16_2_bar CIM_cell
X319 I3163_inv O_3_16_3 WL_3_3 BL BLB W_3_16_3 W_3_16_3_bar CIM_cell
X320 I3164_inv O_3_16_4 WL_3_4 BL BLB W_3_16_4 W_3_16_4_bar CIM_cell
X321 I3171_inv O_3_17_1 WL_3_1 BL BLB W_3_17_1 W_3_17_1_bar CIM_cell
X322 I3172_inv O_3_17_2 WL_3_2 BL BLB W_3_17_2 W_3_17_2_bar CIM_cell
X323 I3173_inv O_3_17_3 WL_3_3 BL BLB W_3_17_3 W_3_17_3_bar CIM_cell
X324 I3174_inv O_3_17_4 WL_3_4 BL BLB W_3_17_4 W_3_17_4_bar CIM_cell
X325 I3181_inv O_3_18_1 WL_3_1 BL BLB W_3_18_1 W_3_18_1_bar CIM_cell
X326 I3182_inv O_3_18_2 WL_3_2 BL BLB W_3_18_2 W_3_18_2_bar CIM_cell
X327 I3183_inv O_3_18_3 WL_3_3 BL BLB W_3_18_3 W_3_18_3_bar CIM_cell
X328 I3184_inv O_3_18_4 WL_3_4 BL BLB W_3_18_4 W_3_18_4_bar CIM_cell
X329 I3191_inv O_3_19_1 WL_3_1 BL BLB W_3_19_1 W_3_19_1_bar CIM_cell
X330 I3192_inv O_3_19_2 WL_3_2 BL BLB W_3_19_2 W_3_19_2_bar CIM_cell
X331 I3193_inv O_3_19_3 WL_3_3 BL BLB W_3_19_3 W_3_19_3_bar CIM_cell
X332 I3194_inv O_3_19_4 WL_3_4 BL BLB W_3_19_4 W_3_19_4_bar CIM_cell
X333 I3201_inv O_3_20_1 WL_3_1 BL BLB W_3_20_1 W_3_20_1_bar CIM_cell
X334 I3202_inv O_3_20_2 WL_3_2 BL BLB W_3_20_2 W_3_20_2_bar CIM_cell
X335 I3203_inv O_3_20_3 WL_3_3 BL BLB W_3_20_3 W_3_20_3_bar CIM_cell
X336 I3204_inv O_3_20_4 WL_3_4 BL BLB W_3_20_4 W_3_20_4_bar CIM_cell
X337 I3211_inv O_3_21_1 WL_3_1 BL BLB W_3_21_1 W_3_21_1_bar CIM_cell
X338 I3212_inv O_3_21_2 WL_3_2 BL BLB W_3_21_2 W_3_21_2_bar CIM_cell
X339 I3213_inv O_3_21_3 WL_3_3 BL BLB W_3_21_3 W_3_21_3_bar CIM_cell
X340 I3214_inv O_3_21_4 WL_3_4 BL BLB W_3_21_4 W_3_21_4_bar CIM_cell
X341 I3221_inv O_3_22_1 WL_3_1 BL BLB W_3_22_1 W_3_22_1_bar CIM_cell
X342 I3222_inv O_3_22_2 WL_3_2 BL BLB W_3_22_2 W_3_22_2_bar CIM_cell
X343 I3223_inv O_3_22_3 WL_3_3 BL BLB W_3_22_3 W_3_22_3_bar CIM_cell
X344 I3224_inv O_3_22_4 WL_3_4 BL BLB W_3_22_4 W_3_22_4_bar CIM_cell
X345 I3231_inv O_3_23_1 WL_3_1 BL BLB W_3_23_1 W_3_23_1_bar CIM_cell
X346 I3232_inv O_3_23_2 WL_3_2 BL BLB W_3_23_2 W_3_23_2_bar CIM_cell
X347 I3233_inv O_3_23_3 WL_3_3 BL BLB W_3_23_3 W_3_23_3_bar CIM_cell
X348 I3234_inv O_3_23_4 WL_3_4 BL BLB W_3_23_4 W_3_23_4_bar CIM_cell
X349 I3241_inv O_3_24_1 WL_3_1 BL BLB W_3_24_1 W_3_24_1_bar CIM_cell
X350 I3242_inv O_3_24_2 WL_3_2 BL BLB W_3_24_2 W_3_24_2_bar CIM_cell
X351 I3243_inv O_3_24_3 WL_3_3 BL BLB W_3_24_3 W_3_24_3_bar CIM_cell
X352 I3244_inv O_3_24_4 WL_3_4 BL BLB W_3_24_4 W_3_24_4_bar CIM_cell
X353 I3251_inv O_3_25_1 WL_3_1 BL BLB W_3_25_1 W_3_25_1_bar CIM_cell
X354 I3252_inv O_3_25_2 WL_3_2 BL BLB W_3_25_2 W_3_25_2_bar CIM_cell
X355 I3253_inv O_3_25_3 WL_3_3 BL BLB W_3_25_3 W_3_25_3_bar CIM_cell
X356 I3254_inv O_3_25_4 WL_3_4 BL BLB W_3_25_4 W_3_25_4_bar CIM_cell
X357 I3261_inv O_3_26_1 WL_3_1 BL BLB W_3_26_1 W_3_26_1_bar CIM_cell
X358 I3262_inv O_3_26_2 WL_3_2 BL BLB W_3_26_2 W_3_26_2_bar CIM_cell
X359 I3263_inv O_3_26_3 WL_3_3 BL BLB W_3_26_3 W_3_26_3_bar CIM_cell
X360 I3264_inv O_3_26_4 WL_3_4 BL BLB W_3_26_4 W_3_26_4_bar CIM_cell
X361 I3271_inv O_3_27_1 WL_3_1 BL BLB W_3_27_1 W_3_27_1_bar CIM_cell
X362 I3272_inv O_3_27_2 WL_3_2 BL BLB W_3_27_2 W_3_27_2_bar CIM_cell
X363 I3273_inv O_3_27_3 WL_3_3 BL BLB W_3_27_3 W_3_27_3_bar CIM_cell
X364 I3274_inv O_3_27_4 WL_3_4 BL BLB W_3_27_4 W_3_27_4_bar CIM_cell
X365 I3281_inv O_3_28_1 WL_3_1 BL BLB W_3_28_1 W_3_28_1_bar CIM_cell
X366 I3282_inv O_3_28_2 WL_3_2 BL BLB W_3_28_2 W_3_28_2_bar CIM_cell
X367 I3283_inv O_3_28_3 WL_3_3 BL BLB W_3_28_3 W_3_28_3_bar CIM_cell
X368 I3284_inv O_3_28_4 WL_3_4 BL BLB W_3_28_4 W_3_28_4_bar CIM_cell
X369 I3291_inv O_3_29_1 WL_3_1 BL BLB W_3_29_1 W_3_29_1_bar CIM_cell
X370 I3292_inv O_3_29_2 WL_3_2 BL BLB W_3_29_2 W_3_29_2_bar CIM_cell
X371 I3293_inv O_3_29_3 WL_3_3 BL BLB W_3_29_3 W_3_29_3_bar CIM_cell
X372 I3294_inv O_3_29_4 WL_3_4 BL BLB W_3_29_4 W_3_29_4_bar CIM_cell
X373 I3301_inv O_3_30_1 WL_3_1 BL BLB W_3_30_1 W_3_30_1_bar CIM_cell
X374 I3302_inv O_3_30_2 WL_3_2 BL BLB W_3_30_2 W_3_30_2_bar CIM_cell
X375 I3303_inv O_3_30_3 WL_3_3 BL BLB W_3_30_3 W_3_30_3_bar CIM_cell
X376 I3304_inv O_3_30_4 WL_3_4 BL BLB W_3_30_4 W_3_30_4_bar CIM_cell
X377 I3311_inv O_3_31_1 WL_3_1 BL BLB W_3_31_1 W_3_31_1_bar CIM_cell
X378 I3312_inv O_3_31_2 WL_3_2 BL BLB W_3_31_2 W_3_31_2_bar CIM_cell
X379 I3313_inv O_3_31_3 WL_3_3 BL BLB W_3_31_3 W_3_31_3_bar CIM_cell
X380 I3314_inv O_3_31_4 WL_3_4 BL BLB W_3_31_4 W_3_31_4_bar CIM_cell
X381 I3321_inv O_3_32_1 WL_3_1 BL BLB W_3_32_1 W_3_32_1_bar CIM_cell
X382 I3322_inv O_3_32_2 WL_3_2 BL BLB W_3_32_2 W_3_32_2_bar CIM_cell
X383 I3323_inv O_3_32_3 WL_3_3 BL BLB W_3_32_3 W_3_32_3_bar CIM_cell
X384 I3324_inv O_3_32_4 WL_3_4 BL BLB W_3_32_4 W_3_32_4_bar CIM_cell
X385 I411_inv O_4_1_1 WL_4_1 BL BLB W_4_1_1 W_4_1_1_bar CIM_cell
X386 I412_inv O_4_1_2 WL_4_2 BL BLB W_4_1_2 W_4_1_2_bar CIM_cell
X387 I413_inv O_4_1_3 WL_4_3 BL BLB W_4_1_3 W_4_1_3_bar CIM_cell
X388 I414_inv O_4_1_4 WL_4_4 BL BLB W_4_1_4 W_4_1_4_bar CIM_cell
X389 I421_inv O_4_2_1 WL_4_1 BL BLB W_4_2_1 W_4_2_1_bar CIM_cell
X390 I422_inv O_4_2_2 WL_4_2 BL BLB W_4_2_2 W_4_2_2_bar CIM_cell
X391 I423_inv O_4_2_3 WL_4_3 BL BLB W_4_2_3 W_4_2_3_bar CIM_cell
X392 I424_inv O_4_2_4 WL_4_4 BL BLB W_4_2_4 W_4_2_4_bar CIM_cell
X393 I431_inv O_4_3_1 WL_4_1 BL BLB W_4_3_1 W_4_3_1_bar CIM_cell
X394 I432_inv O_4_3_2 WL_4_2 BL BLB W_4_3_2 W_4_3_2_bar CIM_cell
X395 I433_inv O_4_3_3 WL_4_3 BL BLB W_4_3_3 W_4_3_3_bar CIM_cell
X396 I434_inv O_4_3_4 WL_4_4 BL BLB W_4_3_4 W_4_3_4_bar CIM_cell
X397 I441_inv O_4_4_1 WL_4_1 BL BLB W_4_4_1 W_4_4_1_bar CIM_cell
X398 I442_inv O_4_4_2 WL_4_2 BL BLB W_4_4_2 W_4_4_2_bar CIM_cell
X399 I443_inv O_4_4_3 WL_4_3 BL BLB W_4_4_3 W_4_4_3_bar CIM_cell
X400 I444_inv O_4_4_4 WL_4_4 BL BLB W_4_4_4 W_4_4_4_bar CIM_cell
X401 I451_inv O_4_5_1 WL_4_1 BL BLB W_4_5_1 W_4_5_1_bar CIM_cell
X402 I452_inv O_4_5_2 WL_4_2 BL BLB W_4_5_2 W_4_5_2_bar CIM_cell
X403 I453_inv O_4_5_3 WL_4_3 BL BLB W_4_5_3 W_4_5_3_bar CIM_cell
X404 I454_inv O_4_5_4 WL_4_4 BL BLB W_4_5_4 W_4_5_4_bar CIM_cell
X405 I461_inv O_4_6_1 WL_4_1 BL BLB W_4_6_1 W_4_6_1_bar CIM_cell
X406 I462_inv O_4_6_2 WL_4_2 BL BLB W_4_6_2 W_4_6_2_bar CIM_cell
X407 I463_inv O_4_6_3 WL_4_3 BL BLB W_4_6_3 W_4_6_3_bar CIM_cell
X408 I464_inv O_4_6_4 WL_4_4 BL BLB W_4_6_4 W_4_6_4_bar CIM_cell
X409 I471_inv O_4_7_1 WL_4_1 BL BLB W_4_7_1 W_4_7_1_bar CIM_cell
X410 I472_inv O_4_7_2 WL_4_2 BL BLB W_4_7_2 W_4_7_2_bar CIM_cell
X411 I473_inv O_4_7_3 WL_4_3 BL BLB W_4_7_3 W_4_7_3_bar CIM_cell
X412 I474_inv O_4_7_4 WL_4_4 BL BLB W_4_7_4 W_4_7_4_bar CIM_cell
X413 I481_inv O_4_8_1 WL_4_1 BL BLB W_4_8_1 W_4_8_1_bar CIM_cell
X414 I482_inv O_4_8_2 WL_4_2 BL BLB W_4_8_2 W_4_8_2_bar CIM_cell
X415 I483_inv O_4_8_3 WL_4_3 BL BLB W_4_8_3 W_4_8_3_bar CIM_cell
X416 I484_inv O_4_8_4 WL_4_4 BL BLB W_4_8_4 W_4_8_4_bar CIM_cell
X417 I491_inv O_4_9_1 WL_4_1 BL BLB W_4_9_1 W_4_9_1_bar CIM_cell
X418 I492_inv O_4_9_2 WL_4_2 BL BLB W_4_9_2 W_4_9_2_bar CIM_cell
X419 I493_inv O_4_9_3 WL_4_3 BL BLB W_4_9_3 W_4_9_3_bar CIM_cell
X420 I494_inv O_4_9_4 WL_4_4 BL BLB W_4_9_4 W_4_9_4_bar CIM_cell
X421 I4101_inv O_4_10_1 WL_4_1 BL BLB W_4_10_1 W_4_10_1_bar CIM_cell
X422 I4102_inv O_4_10_2 WL_4_2 BL BLB W_4_10_2 W_4_10_2_bar CIM_cell
X423 I4103_inv O_4_10_3 WL_4_3 BL BLB W_4_10_3 W_4_10_3_bar CIM_cell
X424 I4104_inv O_4_10_4 WL_4_4 BL BLB W_4_10_4 W_4_10_4_bar CIM_cell
X425 I4111_inv O_4_11_1 WL_4_1 BL BLB W_4_11_1 W_4_11_1_bar CIM_cell
X426 I4112_inv O_4_11_2 WL_4_2 BL BLB W_4_11_2 W_4_11_2_bar CIM_cell
X427 I4113_inv O_4_11_3 WL_4_3 BL BLB W_4_11_3 W_4_11_3_bar CIM_cell
X428 I4114_inv O_4_11_4 WL_4_4 BL BLB W_4_11_4 W_4_11_4_bar CIM_cell
X429 I4121_inv O_4_12_1 WL_4_1 BL BLB W_4_12_1 W_4_12_1_bar CIM_cell
X430 I4122_inv O_4_12_2 WL_4_2 BL BLB W_4_12_2 W_4_12_2_bar CIM_cell
X431 I4123_inv O_4_12_3 WL_4_3 BL BLB W_4_12_3 W_4_12_3_bar CIM_cell
X432 I4124_inv O_4_12_4 WL_4_4 BL BLB W_4_12_4 W_4_12_4_bar CIM_cell
X433 I4131_inv O_4_13_1 WL_4_1 BL BLB W_4_13_1 W_4_13_1_bar CIM_cell
X434 I4132_inv O_4_13_2 WL_4_2 BL BLB W_4_13_2 W_4_13_2_bar CIM_cell
X435 I4133_inv O_4_13_3 WL_4_3 BL BLB W_4_13_3 W_4_13_3_bar CIM_cell
X436 I4134_inv O_4_13_4 WL_4_4 BL BLB W_4_13_4 W_4_13_4_bar CIM_cell
X437 I4141_inv O_4_14_1 WL_4_1 BL BLB W_4_14_1 W_4_14_1_bar CIM_cell
X438 I4142_inv O_4_14_2 WL_4_2 BL BLB W_4_14_2 W_4_14_2_bar CIM_cell
X439 I4143_inv O_4_14_3 WL_4_3 BL BLB W_4_14_3 W_4_14_3_bar CIM_cell
X440 I4144_inv O_4_14_4 WL_4_4 BL BLB W_4_14_4 W_4_14_4_bar CIM_cell
X441 I4151_inv O_4_15_1 WL_4_1 BL BLB W_4_15_1 W_4_15_1_bar CIM_cell
X442 I4152_inv O_4_15_2 WL_4_2 BL BLB W_4_15_2 W_4_15_2_bar CIM_cell
X443 I4153_inv O_4_15_3 WL_4_3 BL BLB W_4_15_3 W_4_15_3_bar CIM_cell
X444 I4154_inv O_4_15_4 WL_4_4 BL BLB W_4_15_4 W_4_15_4_bar CIM_cell
X445 I4161_inv O_4_16_1 WL_4_1 BL BLB W_4_16_1 W_4_16_1_bar CIM_cell
X446 I4162_inv O_4_16_2 WL_4_2 BL BLB W_4_16_2 W_4_16_2_bar CIM_cell
X447 I4163_inv O_4_16_3 WL_4_3 BL BLB W_4_16_3 W_4_16_3_bar CIM_cell
X448 I4164_inv O_4_16_4 WL_4_4 BL BLB W_4_16_4 W_4_16_4_bar CIM_cell
X449 I4171_inv O_4_17_1 WL_4_1 BL BLB W_4_17_1 W_4_17_1_bar CIM_cell
X450 I4172_inv O_4_17_2 WL_4_2 BL BLB W_4_17_2 W_4_17_2_bar CIM_cell
X451 I4173_inv O_4_17_3 WL_4_3 BL BLB W_4_17_3 W_4_17_3_bar CIM_cell
X452 I4174_inv O_4_17_4 WL_4_4 BL BLB W_4_17_4 W_4_17_4_bar CIM_cell
X453 I4181_inv O_4_18_1 WL_4_1 BL BLB W_4_18_1 W_4_18_1_bar CIM_cell
X454 I4182_inv O_4_18_2 WL_4_2 BL BLB W_4_18_2 W_4_18_2_bar CIM_cell
X455 I4183_inv O_4_18_3 WL_4_3 BL BLB W_4_18_3 W_4_18_3_bar CIM_cell
X456 I4184_inv O_4_18_4 WL_4_4 BL BLB W_4_18_4 W_4_18_4_bar CIM_cell
X457 I4191_inv O_4_19_1 WL_4_1 BL BLB W_4_19_1 W_4_19_1_bar CIM_cell
X458 I4192_inv O_4_19_2 WL_4_2 BL BLB W_4_19_2 W_4_19_2_bar CIM_cell
X459 I4193_inv O_4_19_3 WL_4_3 BL BLB W_4_19_3 W_4_19_3_bar CIM_cell
X460 I4194_inv O_4_19_4 WL_4_4 BL BLB W_4_19_4 W_4_19_4_bar CIM_cell
X461 I4201_inv O_4_20_1 WL_4_1 BL BLB W_4_20_1 W_4_20_1_bar CIM_cell
X462 I4202_inv O_4_20_2 WL_4_2 BL BLB W_4_20_2 W_4_20_2_bar CIM_cell
X463 I4203_inv O_4_20_3 WL_4_3 BL BLB W_4_20_3 W_4_20_3_bar CIM_cell
X464 I4204_inv O_4_20_4 WL_4_4 BL BLB W_4_20_4 W_4_20_4_bar CIM_cell
X465 I4211_inv O_4_21_1 WL_4_1 BL BLB W_4_21_1 W_4_21_1_bar CIM_cell
X466 I4212_inv O_4_21_2 WL_4_2 BL BLB W_4_21_2 W_4_21_2_bar CIM_cell
X467 I4213_inv O_4_21_3 WL_4_3 BL BLB W_4_21_3 W_4_21_3_bar CIM_cell
X468 I4214_inv O_4_21_4 WL_4_4 BL BLB W_4_21_4 W_4_21_4_bar CIM_cell
X469 I4221_inv O_4_22_1 WL_4_1 BL BLB W_4_22_1 W_4_22_1_bar CIM_cell
X470 I4222_inv O_4_22_2 WL_4_2 BL BLB W_4_22_2 W_4_22_2_bar CIM_cell
X471 I4223_inv O_4_22_3 WL_4_3 BL BLB W_4_22_3 W_4_22_3_bar CIM_cell
X472 I4224_inv O_4_22_4 WL_4_4 BL BLB W_4_22_4 W_4_22_4_bar CIM_cell
X473 I4231_inv O_4_23_1 WL_4_1 BL BLB W_4_23_1 W_4_23_1_bar CIM_cell
X474 I4232_inv O_4_23_2 WL_4_2 BL BLB W_4_23_2 W_4_23_2_bar CIM_cell
X475 I4233_inv O_4_23_3 WL_4_3 BL BLB W_4_23_3 W_4_23_3_bar CIM_cell
X476 I4234_inv O_4_23_4 WL_4_4 BL BLB W_4_23_4 W_4_23_4_bar CIM_cell
X477 I4241_inv O_4_24_1 WL_4_1 BL BLB W_4_24_1 W_4_24_1_bar CIM_cell
X478 I4242_inv O_4_24_2 WL_4_2 BL BLB W_4_24_2 W_4_24_2_bar CIM_cell
X479 I4243_inv O_4_24_3 WL_4_3 BL BLB W_4_24_3 W_4_24_3_bar CIM_cell
X480 I4244_inv O_4_24_4 WL_4_4 BL BLB W_4_24_4 W_4_24_4_bar CIM_cell
X481 I4251_inv O_4_25_1 WL_4_1 BL BLB W_4_25_1 W_4_25_1_bar CIM_cell
X482 I4252_inv O_4_25_2 WL_4_2 BL BLB W_4_25_2 W_4_25_2_bar CIM_cell
X483 I4253_inv O_4_25_3 WL_4_3 BL BLB W_4_25_3 W_4_25_3_bar CIM_cell
X484 I4254_inv O_4_25_4 WL_4_4 BL BLB W_4_25_4 W_4_25_4_bar CIM_cell
X485 I4261_inv O_4_26_1 WL_4_1 BL BLB W_4_26_1 W_4_26_1_bar CIM_cell
X486 I4262_inv O_4_26_2 WL_4_2 BL BLB W_4_26_2 W_4_26_2_bar CIM_cell
X487 I4263_inv O_4_26_3 WL_4_3 BL BLB W_4_26_3 W_4_26_3_bar CIM_cell
X488 I4264_inv O_4_26_4 WL_4_4 BL BLB W_4_26_4 W_4_26_4_bar CIM_cell
X489 I4271_inv O_4_27_1 WL_4_1 BL BLB W_4_27_1 W_4_27_1_bar CIM_cell
X490 I4272_inv O_4_27_2 WL_4_2 BL BLB W_4_27_2 W_4_27_2_bar CIM_cell
X491 I4273_inv O_4_27_3 WL_4_3 BL BLB W_4_27_3 W_4_27_3_bar CIM_cell
X492 I4274_inv O_4_27_4 WL_4_4 BL BLB W_4_27_4 W_4_27_4_bar CIM_cell
X493 I4281_inv O_4_28_1 WL_4_1 BL BLB W_4_28_1 W_4_28_1_bar CIM_cell
X494 I4282_inv O_4_28_2 WL_4_2 BL BLB W_4_28_2 W_4_28_2_bar CIM_cell
X495 I4283_inv O_4_28_3 WL_4_3 BL BLB W_4_28_3 W_4_28_3_bar CIM_cell
X496 I4284_inv O_4_28_4 WL_4_4 BL BLB W_4_28_4 W_4_28_4_bar CIM_cell
X497 I4291_inv O_4_29_1 WL_4_1 BL BLB W_4_29_1 W_4_29_1_bar CIM_cell
X498 I4292_inv O_4_29_2 WL_4_2 BL BLB W_4_29_2 W_4_29_2_bar CIM_cell
X499 I4293_inv O_4_29_3 WL_4_3 BL BLB W_4_29_3 W_4_29_3_bar CIM_cell
X500 I4294_inv O_4_29_4 WL_4_4 BL BLB W_4_29_4 W_4_29_4_bar CIM_cell
X501 I4301_inv O_4_30_1 WL_4_1 BL BLB W_4_30_1 W_4_30_1_bar CIM_cell
X502 I4302_inv O_4_30_2 WL_4_2 BL BLB W_4_30_2 W_4_30_2_bar CIM_cell
X503 I4303_inv O_4_30_3 WL_4_3 BL BLB W_4_30_3 W_4_30_3_bar CIM_cell
X504 I4304_inv O_4_30_4 WL_4_4 BL BLB W_4_30_4 W_4_30_4_bar CIM_cell
X505 I4311_inv O_4_31_1 WL_4_1 BL BLB W_4_31_1 W_4_31_1_bar CIM_cell
X506 I4312_inv O_4_31_2 WL_4_2 BL BLB W_4_31_2 W_4_31_2_bar CIM_cell
X507 I4313_inv O_4_31_3 WL_4_3 BL BLB W_4_31_3 W_4_31_3_bar CIM_cell
X508 I4314_inv O_4_31_4 WL_4_4 BL BLB W_4_31_4 W_4_31_4_bar CIM_cell
X509 I4321_inv O_4_32_1 WL_4_1 BL BLB W_4_32_1 W_4_32_1_bar CIM_cell
X510 I4322_inv O_4_32_2 WL_4_2 BL BLB W_4_32_2 W_4_32_2_bar CIM_cell
X511 I4323_inv O_4_32_3 WL_4_3 BL BLB W_4_32_3 W_4_32_3_bar CIM_cell
X512 I4324_inv O_4_32_4 WL_4_4 BL BLB W_4_32_4 W_4_32_4_bar CIM_cell






***-----------------------***
***      sub-circuit      ***
***-----------------------***

* // QB : weight 
* // input 
* // output 
* .subckt CIM_cell Input Output WL BL BLB q qb
*     X01 WL BL BLB q qb SRAM_6T
*     X02 qb Input Output NOR_2
* .ends

.subckt CIM_cell Input Output WL BL BLB q qb
    X01 WL BL BLB q qb SRAM_6T
    X02 qb Input Output NOR_2
.ends


.subckt SRAM_6T WL BL BLB q qb
    MP1 q   qb  VDD VDD pmos_sram m=1
    MP2 qb  q   VDD VDD pmos_sram m=1
    MN1 q   qb  GND GND nmos_sram m=1
    MN2 qb  q   GND GND nmos_sram m=1
    MN3 BL  WL  q   GND nmos_sram m=1
    MN4 qb  WL  BLB GND nmos_sram m=1
.ends

.subckt NOR_2 A B Y
    MP1 N1  A   VDD VDD pmos_lvt m=1
    MP2 Y   B   N1  VDD pmos_lvt m=1
    MN1 Y   A   GND GND nmos_lvt m=1
    MN2 Y   B   GND GND nmos_lvt m=1
.ends

.subckt Buffer in out
    X_INV1 in   in_b INV
    X_INV2 in_b out  INV
.ends

.subckt INV in out
    Mp  out  in  VDD  VDD  pmos_lvt  m=1
    Mn  out  in  GND  GND  nmos_lvt  m=1
.ends

* Example .IC file for initializing SRAM weights
.IC V(W_1_1_1) = 0 V(W_1_1_1_bar) = 1
.IC V(W_1_1_2) = 1 V(W_1_1_2_bar) = 0
.IC V(W_1_1_3) = 0 V(W_1_1_3_bar) = 1
.IC V(W_1_1_4) = 1 V(W_1_1_4_bar) = 0
.IC V(W_1_2_1) = 0 V(W_1_2_1_bar) = 1
.IC V(W_1_2_2) = 1 V(W_1_2_2_bar) = 0
.IC V(W_1_2_3) = 0 V(W_1_2_3_bar) = 1
.IC V(W_1_2_4) = 1 V(W_1_2_4_bar) = 0
.IC V(W_1_3_1) = 0 V(W_1_3_1_bar) = 1
.IC V(W_1_3_2) = 1 V(W_1_3_2_bar) = 0
.IC V(W_1_3_3) = 0 V(W_1_3_3_bar) = 1
.IC V(W_1_3_4) = 1 V(W_1_3_4_bar) = 0
.IC V(W_1_4_1) = 0 V(W_1_4_1_bar) = 1
.IC V(W_1_4_2) = 1 V(W_1_4_2_bar) = 0
.IC V(W_1_4_3) = 0 V(W_1_4_3_bar) = 1
.IC V(W_1_4_4) = 1 V(W_1_4_4_bar) = 0
.IC V(W_1_5_1) = 0 V(W_1_5_1_bar) = 1
.IC V(W_1_5_2) = 1 V(W_1_5_2_bar) = 0
.IC V(W_1_5_3) = 0 V(W_1_5_3_bar) = 1
.IC V(W_1_5_4) = 1 V(W_1_5_4_bar) = 0
.IC V(W_1_6_1) = 0 V(W_1_6_1_bar) = 1
.IC V(W_1_6_2) = 1 V(W_1_6_2_bar) = 0
.IC V(W_1_6_3) = 0 V(W_1_6_3_bar) = 1
.IC V(W_1_6_4) = 1 V(W_1_6_4_bar) = 0
.IC V(W_1_7_1) = 0 V(W_1_7_1_bar) = 1
.IC V(W_1_7_2) = 1 V(W_1_7_2_bar) = 0
.IC V(W_1_7_3) = 0 V(W_1_7_3_bar) = 1
.IC V(W_1_7_4) = 1 V(W_1_7_4_bar) = 0
.IC V(W_1_8_1) = 0 V(W_1_8_1_bar) = 1
.IC V(W_1_8_2) = 1 V(W_1_8_2_bar) = 0
.IC V(W_1_8_3) = 0 V(W_1_8_3_bar) = 1
.IC V(W_1_8_4) = 1 V(W_1_8_4_bar) = 0
.IC V(W_1_9_1) = 0 V(W_1_9_1_bar) = 1
.IC V(W_1_9_2) = 1 V(W_1_9_2_bar) = 0
.IC V(W_1_9_3) = 0 V(W_1_9_3_bar) = 1
.IC V(W_1_9_4) = 1 V(W_1_9_4_bar) = 0
.IC V(W_1_10_1) = 0 V(W_1_10_1_bar) = 1
.IC V(W_1_10_2) = 1 V(W_1_10_2_bar) = 0
.IC V(W_1_10_3) = 0 V(W_1_10_3_bar) = 1
.IC V(W_1_10_4) = 1 V(W_1_10_4_bar) = 0
.IC V(W_1_11_1) = 0 V(W_1_11_1_bar) = 1
.IC V(W_1_11_2) = 1 V(W_1_11_2_bar) = 0
.IC V(W_1_11_3) = 0 V(W_1_11_3_bar) = 1
.IC V(W_1_11_4) = 1 V(W_1_11_4_bar) = 0
.IC V(W_1_12_1) = 0 V(W_1_12_1_bar) = 1
.IC V(W_1_12_2) = 1 V(W_1_12_2_bar) = 0
.IC V(W_1_12_3) = 0 V(W_1_12_3_bar) = 1
.IC V(W_1_12_4) = 1 V(W_1_12_4_bar) = 0
.IC V(W_1_13_1) = 0 V(W_1_13_1_bar) = 1
.IC V(W_1_13_2) = 1 V(W_1_13_2_bar) = 0
.IC V(W_1_13_3) = 0 V(W_1_13_3_bar) = 1
.IC V(W_1_13_4) = 1 V(W_1_13_4_bar) = 0
.IC V(W_1_14_1) = 0 V(W_1_14_1_bar) = 1
.IC V(W_1_14_2) = 1 V(W_1_14_2_bar) = 0
.IC V(W_1_14_3) = 0 V(W_1_14_3_bar) = 1
.IC V(W_1_14_4) = 1 V(W_1_14_4_bar) = 0
.IC V(W_1_15_1) = 0 V(W_1_15_1_bar) = 1
.IC V(W_1_15_2) = 1 V(W_1_15_2_bar) = 0
.IC V(W_1_15_3) = 0 V(W_1_15_3_bar) = 1
.IC V(W_1_15_4) = 1 V(W_1_15_4_bar) = 0
.IC V(W_1_16_1) = 0 V(W_1_16_1_bar) = 1
.IC V(W_1_16_2) = 1 V(W_1_16_2_bar) = 0
.IC V(W_1_16_3) = 0 V(W_1_16_3_bar) = 1
.IC V(W_1_16_4) = 1 V(W_1_16_4_bar) = 0
.IC V(W_1_17_1) = 0 V(W_1_17_1_bar) = 1
.IC V(W_1_17_2) = 1 V(W_1_17_2_bar) = 0
.IC V(W_1_17_3) = 0 V(W_1_17_3_bar) = 1
.IC V(W_1_17_4) = 1 V(W_1_17_4_bar) = 0
.IC V(W_1_18_1) = 0 V(W_1_18_1_bar) = 1
.IC V(W_1_18_2) = 1 V(W_1_18_2_bar) = 0
.IC V(W_1_18_3) = 0 V(W_1_18_3_bar) = 1
.IC V(W_1_18_4) = 1 V(W_1_18_4_bar) = 0
.IC V(W_1_19_1) = 0 V(W_1_19_1_bar) = 1
.IC V(W_1_19_2) = 1 V(W_1_19_2_bar) = 0
.IC V(W_1_19_3) = 0 V(W_1_19_3_bar) = 1
.IC V(W_1_19_4) = 1 V(W_1_19_4_bar) = 0
.IC V(W_1_20_1) = 0 V(W_1_20_1_bar) = 1
.IC V(W_1_20_2) = 1 V(W_1_20_2_bar) = 0
.IC V(W_1_20_3) = 0 V(W_1_20_3_bar) = 1
.IC V(W_1_20_4) = 1 V(W_1_20_4_bar) = 0
.IC V(W_1_21_1) = 0 V(W_1_21_1_bar) = 1
.IC V(W_1_21_2) = 1 V(W_1_21_2_bar) = 0
.IC V(W_1_21_3) = 0 V(W_1_21_3_bar) = 1
.IC V(W_1_21_4) = 1 V(W_1_21_4_bar) = 0
.IC V(W_1_22_1) = 0 V(W_1_22_1_bar) = 1
.IC V(W_1_22_2) = 1 V(W_1_22_2_bar) = 0
.IC V(W_1_22_3) = 0 V(W_1_22_3_bar) = 1
.IC V(W_1_22_4) = 1 V(W_1_22_4_bar) = 0
.IC V(W_1_23_1) = 0 V(W_1_23_1_bar) = 1
.IC V(W_1_23_2) = 1 V(W_1_23_2_bar) = 0
.IC V(W_1_23_3) = 0 V(W_1_23_3_bar) = 1
.IC V(W_1_23_4) = 1 V(W_1_23_4_bar) = 0
.IC V(W_1_24_1) = 0 V(W_1_24_1_bar) = 1
.IC V(W_1_24_2) = 1 V(W_1_24_2_bar) = 0
.IC V(W_1_24_3) = 0 V(W_1_24_3_bar) = 1
.IC V(W_1_24_4) = 1 V(W_1_24_4_bar) = 0
.IC V(W_1_25_1) = 0 V(W_1_25_1_bar) = 1
.IC V(W_1_25_2) = 1 V(W_1_25_2_bar) = 0
.IC V(W_1_25_3) = 0 V(W_1_25_3_bar) = 1
.IC V(W_1_25_4) = 1 V(W_1_25_4_bar) = 0
.IC V(W_1_26_1) = 0 V(W_1_26_1_bar) = 1
.IC V(W_1_26_2) = 1 V(W_1_26_2_bar) = 0
.IC V(W_1_26_3) = 0 V(W_1_26_3_bar) = 1
.IC V(W_1_26_4) = 1 V(W_1_26_4_bar) = 0
.IC V(W_1_27_1) = 0 V(W_1_27_1_bar) = 1
.IC V(W_1_27_2) = 1 V(W_1_27_2_bar) = 0
.IC V(W_1_27_3) = 0 V(W_1_27_3_bar) = 1
.IC V(W_1_27_4) = 1 V(W_1_27_4_bar) = 0
.IC V(W_1_28_1) = 0 V(W_1_28_1_bar) = 1
.IC V(W_1_28_2) = 1 V(W_1_28_2_bar) = 0
.IC V(W_1_28_3) = 0 V(W_1_28_3_bar) = 1
.IC V(W_1_28_4) = 1 V(W_1_28_4_bar) = 0
.IC V(W_1_29_1) = 0 V(W_1_29_1_bar) = 1
.IC V(W_1_29_2) = 1 V(W_1_29_2_bar) = 0
.IC V(W_1_29_3) = 0 V(W_1_29_3_bar) = 1
.IC V(W_1_29_4) = 1 V(W_1_29_4_bar) = 0
.IC V(W_1_30_1) = 0 V(W_1_30_1_bar) = 1
.IC V(W_1_30_2) = 1 V(W_1_30_2_bar) = 0
.IC V(W_1_30_3) = 0 V(W_1_30_3_bar) = 1
.IC V(W_1_30_4) = 1 V(W_1_30_4_bar) = 0
.IC V(W_1_31_1) = 0 V(W_1_31_1_bar) = 1
.IC V(W_1_31_2) = 1 V(W_1_31_2_bar) = 0
.IC V(W_1_31_3) = 0 V(W_1_31_3_bar) = 1
.IC V(W_1_31_4) = 1 V(W_1_31_4_bar) = 0
.IC V(W_1_32_1) = 0 V(W_1_32_1_bar) = 1
.IC V(W_1_32_2) = 1 V(W_1_32_2_bar) = 0
.IC V(W_1_32_3) = 0 V(W_1_32_3_bar) = 1
.IC V(W_1_32_4) = 1 V(W_1_32_4_bar) = 0
.IC V(W_2_1_1) = 0 V(W_2_1_1_bar) = 1
.IC V(W_2_1_2) = 1 V(W_2_1_2_bar) = 0
.IC V(W_2_1_3) = 0 V(W_2_1_3_bar) = 1
.IC V(W_2_1_4) = 1 V(W_2_1_4_bar) = 0
.IC V(W_2_2_1) = 0 V(W_2_2_1_bar) = 1
.IC V(W_2_2_2) = 1 V(W_2_2_2_bar) = 0
.IC V(W_2_2_3) = 0 V(W_2_2_3_bar) = 1
.IC V(W_2_2_4) = 1 V(W_2_2_4_bar) = 0
.IC V(W_2_3_1) = 0 V(W_2_3_1_bar) = 1
.IC V(W_2_3_2) = 1 V(W_2_3_2_bar) = 0
.IC V(W_2_3_3) = 0 V(W_2_3_3_bar) = 1
.IC V(W_2_3_4) = 1 V(W_2_3_4_bar) = 0
.IC V(W_2_4_1) = 0 V(W_2_4_1_bar) = 1
.IC V(W_2_4_2) = 1 V(W_2_4_2_bar) = 0
.IC V(W_2_4_3) = 0 V(W_2_4_3_bar) = 1
.IC V(W_2_4_4) = 1 V(W_2_4_4_bar) = 0
.IC V(W_2_5_1) = 0 V(W_2_5_1_bar) = 1
.IC V(W_2_5_2) = 1 V(W_2_5_2_bar) = 0
.IC V(W_2_5_3) = 0 V(W_2_5_3_bar) = 1
.IC V(W_2_5_4) = 1 V(W_2_5_4_bar) = 0
.IC V(W_2_6_1) = 0 V(W_2_6_1_bar) = 1
.IC V(W_2_6_2) = 1 V(W_2_6_2_bar) = 0
.IC V(W_2_6_3) = 0 V(W_2_6_3_bar) = 1
.IC V(W_2_6_4) = 1 V(W_2_6_4_bar) = 0
.IC V(W_2_7_1) = 0 V(W_2_7_1_bar) = 1
.IC V(W_2_7_2) = 1 V(W_2_7_2_bar) = 0
.IC V(W_2_7_3) = 0 V(W_2_7_3_bar) = 1
.IC V(W_2_7_4) = 1 V(W_2_7_4_bar) = 0
.IC V(W_2_8_1) = 0 V(W_2_8_1_bar) = 1
.IC V(W_2_8_2) = 1 V(W_2_8_2_bar) = 0
.IC V(W_2_8_3) = 0 V(W_2_8_3_bar) = 1
.IC V(W_2_8_4) = 1 V(W_2_8_4_bar) = 0
.IC V(W_2_9_1) = 0 V(W_2_9_1_bar) = 1
.IC V(W_2_9_2) = 1 V(W_2_9_2_bar) = 0
.IC V(W_2_9_3) = 0 V(W_2_9_3_bar) = 1
.IC V(W_2_9_4) = 1 V(W_2_9_4_bar) = 0
.IC V(W_2_10_1) = 0 V(W_2_10_1_bar) = 1
.IC V(W_2_10_2) = 1 V(W_2_10_2_bar) = 0
.IC V(W_2_10_3) = 0 V(W_2_10_3_bar) = 1
.IC V(W_2_10_4) = 1 V(W_2_10_4_bar) = 0
.IC V(W_2_11_1) = 0 V(W_2_11_1_bar) = 1
.IC V(W_2_11_2) = 1 V(W_2_11_2_bar) = 0
.IC V(W_2_11_3) = 0 V(W_2_11_3_bar) = 1
.IC V(W_2_11_4) = 1 V(W_2_11_4_bar) = 0
.IC V(W_2_12_1) = 0 V(W_2_12_1_bar) = 1
.IC V(W_2_12_2) = 1 V(W_2_12_2_bar) = 0
.IC V(W_2_12_3) = 0 V(W_2_12_3_bar) = 1
.IC V(W_2_12_4) = 1 V(W_2_12_4_bar) = 0
.IC V(W_2_13_1) = 0 V(W_2_13_1_bar) = 1
.IC V(W_2_13_2) = 1 V(W_2_13_2_bar) = 0
.IC V(W_2_13_3) = 0 V(W_2_13_3_bar) = 1
.IC V(W_2_13_4) = 1 V(W_2_13_4_bar) = 0
.IC V(W_2_14_1) = 0 V(W_2_14_1_bar) = 1
.IC V(W_2_14_2) = 1 V(W_2_14_2_bar) = 0
.IC V(W_2_14_3) = 0 V(W_2_14_3_bar) = 1
.IC V(W_2_14_4) = 1 V(W_2_14_4_bar) = 0
.IC V(W_2_15_1) = 0 V(W_2_15_1_bar) = 1
.IC V(W_2_15_2) = 1 V(W_2_15_2_bar) = 0
.IC V(W_2_15_3) = 0 V(W_2_15_3_bar) = 1
.IC V(W_2_15_4) = 1 V(W_2_15_4_bar) = 0
.IC V(W_2_16_1) = 0 V(W_2_16_1_bar) = 1
.IC V(W_2_16_2) = 1 V(W_2_16_2_bar) = 0
.IC V(W_2_16_3) = 0 V(W_2_16_3_bar) = 1
.IC V(W_2_16_4) = 1 V(W_2_16_4_bar) = 0
.IC V(W_2_17_1) = 0 V(W_2_17_1_bar) = 1
.IC V(W_2_17_2) = 1 V(W_2_17_2_bar) = 0
.IC V(W_2_17_3) = 0 V(W_2_17_3_bar) = 1
.IC V(W_2_17_4) = 1 V(W_2_17_4_bar) = 0
.IC V(W_2_18_1) = 0 V(W_2_18_1_bar) = 1
.IC V(W_2_18_2) = 1 V(W_2_18_2_bar) = 0
.IC V(W_2_18_3) = 0 V(W_2_18_3_bar) = 1
.IC V(W_2_18_4) = 1 V(W_2_18_4_bar) = 0
.IC V(W_2_19_1) = 0 V(W_2_19_1_bar) = 1
.IC V(W_2_19_2) = 1 V(W_2_19_2_bar) = 0
.IC V(W_2_19_3) = 0 V(W_2_19_3_bar) = 1
.IC V(W_2_19_4) = 1 V(W_2_19_4_bar) = 0
.IC V(W_2_20_1) = 0 V(W_2_20_1_bar) = 1
.IC V(W_2_20_2) = 1 V(W_2_20_2_bar) = 0
.IC V(W_2_20_3) = 0 V(W_2_20_3_bar) = 1
.IC V(W_2_20_4) = 1 V(W_2_20_4_bar) = 0
.IC V(W_2_21_1) = 0 V(W_2_21_1_bar) = 1
.IC V(W_2_21_2) = 1 V(W_2_21_2_bar) = 0
.IC V(W_2_21_3) = 0 V(W_2_21_3_bar) = 1
.IC V(W_2_21_4) = 1 V(W_2_21_4_bar) = 0
.IC V(W_2_22_1) = 0 V(W_2_22_1_bar) = 1
.IC V(W_2_22_2) = 1 V(W_2_22_2_bar) = 0
.IC V(W_2_22_3) = 0 V(W_2_22_3_bar) = 1
.IC V(W_2_22_4) = 1 V(W_2_22_4_bar) = 0
.IC V(W_2_23_1) = 0 V(W_2_23_1_bar) = 1
.IC V(W_2_23_2) = 1 V(W_2_23_2_bar) = 0
.IC V(W_2_23_3) = 0 V(W_2_23_3_bar) = 1
.IC V(W_2_23_4) = 1 V(W_2_23_4_bar) = 0
.IC V(W_2_24_1) = 0 V(W_2_24_1_bar) = 1
.IC V(W_2_24_2) = 1 V(W_2_24_2_bar) = 0
.IC V(W_2_24_3) = 0 V(W_2_24_3_bar) = 1
.IC V(W_2_24_4) = 1 V(W_2_24_4_bar) = 0
.IC V(W_2_25_1) = 0 V(W_2_25_1_bar) = 1
.IC V(W_2_25_2) = 1 V(W_2_25_2_bar) = 0
.IC V(W_2_25_3) = 0 V(W_2_25_3_bar) = 1
.IC V(W_2_25_4) = 1 V(W_2_25_4_bar) = 0
.IC V(W_2_26_1) = 0 V(W_2_26_1_bar) = 1
.IC V(W_2_26_2) = 1 V(W_2_26_2_bar) = 0
.IC V(W_2_26_3) = 0 V(W_2_26_3_bar) = 1
.IC V(W_2_26_4) = 1 V(W_2_26_4_bar) = 0
.IC V(W_2_27_1) = 0 V(W_2_27_1_bar) = 1
.IC V(W_2_27_2) = 1 V(W_2_27_2_bar) = 0
.IC V(W_2_27_3) = 0 V(W_2_27_3_bar) = 1
.IC V(W_2_27_4) = 1 V(W_2_27_4_bar) = 0
.IC V(W_2_28_1) = 0 V(W_2_28_1_bar) = 1
.IC V(W_2_28_2) = 1 V(W_2_28_2_bar) = 0
.IC V(W_2_28_3) = 0 V(W_2_28_3_bar) = 1
.IC V(W_2_28_4) = 1 V(W_2_28_4_bar) = 0
.IC V(W_2_29_1) = 0 V(W_2_29_1_bar) = 1
.IC V(W_2_29_2) = 1 V(W_2_29_2_bar) = 0
.IC V(W_2_29_3) = 0 V(W_2_29_3_bar) = 1
.IC V(W_2_29_4) = 1 V(W_2_29_4_bar) = 0
.IC V(W_2_30_1) = 0 V(W_2_30_1_bar) = 1
.IC V(W_2_30_2) = 1 V(W_2_30_2_bar) = 0
.IC V(W_2_30_3) = 0 V(W_2_30_3_bar) = 1
.IC V(W_2_30_4) = 1 V(W_2_30_4_bar) = 0
.IC V(W_2_31_1) = 0 V(W_2_31_1_bar) = 1
.IC V(W_2_31_2) = 1 V(W_2_31_2_bar) = 0
.IC V(W_2_31_3) = 0 V(W_2_31_3_bar) = 1
.IC V(W_2_31_4) = 1 V(W_2_31_4_bar) = 0
.IC V(W_2_32_1) = 0 V(W_2_32_1_bar) = 1
.IC V(W_2_32_2) = 1 V(W_2_32_2_bar) = 0
.IC V(W_2_32_3) = 0 V(W_2_32_3_bar) = 1
.IC V(W_2_32_4) = 1 V(W_2_32_4_bar) = 0
.IC V(W_3_1_1) = 0 V(W_3_1_1_bar) = 1
.IC V(W_3_1_2) = 1 V(W_3_1_2_bar) = 0
.IC V(W_3_1_3) = 0 V(W_3_1_3_bar) = 1
.IC V(W_3_1_4) = 1 V(W_3_1_4_bar) = 0
.IC V(W_3_2_1) = 0 V(W_3_2_1_bar) = 1
.IC V(W_3_2_2) = 1 V(W_3_2_2_bar) = 0
.IC V(W_3_2_3) = 0 V(W_3_2_3_bar) = 1
.IC V(W_3_2_4) = 1 V(W_3_2_4_bar) = 0
.IC V(W_3_3_1) = 0 V(W_3_3_1_bar) = 1
.IC V(W_3_3_2) = 1 V(W_3_3_2_bar) = 0
.IC V(W_3_3_3) = 0 V(W_3_3_3_bar) = 1
.IC V(W_3_3_4) = 1 V(W_3_3_4_bar) = 0
.IC V(W_3_4_1) = 0 V(W_3_4_1_bar) = 1
.IC V(W_3_4_2) = 1 V(W_3_4_2_bar) = 0
.IC V(W_3_4_3) = 0 V(W_3_4_3_bar) = 1
.IC V(W_3_4_4) = 1 V(W_3_4_4_bar) = 0
.IC V(W_3_5_1) = 0 V(W_3_5_1_bar) = 1
.IC V(W_3_5_2) = 1 V(W_3_5_2_bar) = 0
.IC V(W_3_5_3) = 0 V(W_3_5_3_bar) = 1
.IC V(W_3_5_4) = 1 V(W_3_5_4_bar) = 0
.IC V(W_3_6_1) = 0 V(W_3_6_1_bar) = 1
.IC V(W_3_6_2) = 1 V(W_3_6_2_bar) = 0
.IC V(W_3_6_3) = 0 V(W_3_6_3_bar) = 1
.IC V(W_3_6_4) = 1 V(W_3_6_4_bar) = 0
.IC V(W_3_7_1) = 0 V(W_3_7_1_bar) = 1
.IC V(W_3_7_2) = 1 V(W_3_7_2_bar) = 0
.IC V(W_3_7_3) = 0 V(W_3_7_3_bar) = 1
.IC V(W_3_7_4) = 1 V(W_3_7_4_bar) = 0
.IC V(W_3_8_1) = 0 V(W_3_8_1_bar) = 1
.IC V(W_3_8_2) = 1 V(W_3_8_2_bar) = 0
.IC V(W_3_8_3) = 0 V(W_3_8_3_bar) = 1
.IC V(W_3_8_4) = 1 V(W_3_8_4_bar) = 0
.IC V(W_3_9_1) = 0 V(W_3_9_1_bar) = 1
.IC V(W_3_9_2) = 1 V(W_3_9_2_bar) = 0
.IC V(W_3_9_3) = 0 V(W_3_9_3_bar) = 1
.IC V(W_3_9_4) = 1 V(W_3_9_4_bar) = 0
.IC V(W_3_10_1) = 0 V(W_3_10_1_bar) = 1
.IC V(W_3_10_2) = 1 V(W_3_10_2_bar) = 0
.IC V(W_3_10_3) = 0 V(W_3_10_3_bar) = 1
.IC V(W_3_10_4) = 1 V(W_3_10_4_bar) = 0
.IC V(W_3_11_1) = 0 V(W_3_11_1_bar) = 1
.IC V(W_3_11_2) = 1 V(W_3_11_2_bar) = 0
.IC V(W_3_11_3) = 0 V(W_3_11_3_bar) = 1
.IC V(W_3_11_4) = 1 V(W_3_11_4_bar) = 0
.IC V(W_3_12_1) = 0 V(W_3_12_1_bar) = 1
.IC V(W_3_12_2) = 1 V(W_3_12_2_bar) = 0
.IC V(W_3_12_3) = 0 V(W_3_12_3_bar) = 1
.IC V(W_3_12_4) = 1 V(W_3_12_4_bar) = 0
.IC V(W_3_13_1) = 0 V(W_3_13_1_bar) = 1
.IC V(W_3_13_2) = 1 V(W_3_13_2_bar) = 0
.IC V(W_3_13_3) = 0 V(W_3_13_3_bar) = 1
.IC V(W_3_13_4) = 1 V(W_3_13_4_bar) = 0
.IC V(W_3_14_1) = 0 V(W_3_14_1_bar) = 1
.IC V(W_3_14_2) = 1 V(W_3_14_2_bar) = 0
.IC V(W_3_14_3) = 0 V(W_3_14_3_bar) = 1
.IC V(W_3_14_4) = 1 V(W_3_14_4_bar) = 0
.IC V(W_3_15_1) = 0 V(W_3_15_1_bar) = 1
.IC V(W_3_15_2) = 1 V(W_3_15_2_bar) = 0
.IC V(W_3_15_3) = 0 V(W_3_15_3_bar) = 1
.IC V(W_3_15_4) = 1 V(W_3_15_4_bar) = 0
.IC V(W_3_16_1) = 0 V(W_3_16_1_bar) = 1
.IC V(W_3_16_2) = 1 V(W_3_16_2_bar) = 0
.IC V(W_3_16_3) = 0 V(W_3_16_3_bar) = 1
.IC V(W_3_16_4) = 1 V(W_3_16_4_bar) = 0
.IC V(W_3_17_1) = 0 V(W_3_17_1_bar) = 1
.IC V(W_3_17_2) = 1 V(W_3_17_2_bar) = 0
.IC V(W_3_17_3) = 0 V(W_3_17_3_bar) = 1
.IC V(W_3_17_4) = 1 V(W_3_17_4_bar) = 0
.IC V(W_3_18_1) = 0 V(W_3_18_1_bar) = 1
.IC V(W_3_18_2) = 1 V(W_3_18_2_bar) = 0
.IC V(W_3_18_3) = 0 V(W_3_18_3_bar) = 1
.IC V(W_3_18_4) = 1 V(W_3_18_4_bar) = 0
.IC V(W_3_19_1) = 0 V(W_3_19_1_bar) = 1
.IC V(W_3_19_2) = 1 V(W_3_19_2_bar) = 0
.IC V(W_3_19_3) = 0 V(W_3_19_3_bar) = 1
.IC V(W_3_19_4) = 1 V(W_3_19_4_bar) = 0
.IC V(W_3_20_1) = 0 V(W_3_20_1_bar) = 1
.IC V(W_3_20_2) = 1 V(W_3_20_2_bar) = 0
.IC V(W_3_20_3) = 0 V(W_3_20_3_bar) = 1
.IC V(W_3_20_4) = 1 V(W_3_20_4_bar) = 0
.IC V(W_3_21_1) = 0 V(W_3_21_1_bar) = 1
.IC V(W_3_21_2) = 1 V(W_3_21_2_bar) = 0
.IC V(W_3_21_3) = 0 V(W_3_21_3_bar) = 1
.IC V(W_3_21_4) = 1 V(W_3_21_4_bar) = 0
.IC V(W_3_22_1) = 0 V(W_3_22_1_bar) = 1
.IC V(W_3_22_2) = 1 V(W_3_22_2_bar) = 0
.IC V(W_3_22_3) = 0 V(W_3_22_3_bar) = 1
.IC V(W_3_22_4) = 1 V(W_3_22_4_bar) = 0
.IC V(W_3_23_1) = 0 V(W_3_23_1_bar) = 1
.IC V(W_3_23_2) = 1 V(W_3_23_2_bar) = 0
.IC V(W_3_23_3) = 0 V(W_3_23_3_bar) = 1
.IC V(W_3_23_4) = 1 V(W_3_23_4_bar) = 0
.IC V(W_3_24_1) = 0 V(W_3_24_1_bar) = 1
.IC V(W_3_24_2) = 1 V(W_3_24_2_bar) = 0
.IC V(W_3_24_3) = 0 V(W_3_24_3_bar) = 1
.IC V(W_3_24_4) = 1 V(W_3_24_4_bar) = 0
.IC V(W_3_25_1) = 0 V(W_3_25_1_bar) = 1
.IC V(W_3_25_2) = 1 V(W_3_25_2_bar) = 0
.IC V(W_3_25_3) = 0 V(W_3_25_3_bar) = 1
.IC V(W_3_25_4) = 1 V(W_3_25_4_bar) = 0
.IC V(W_3_26_1) = 0 V(W_3_26_1_bar) = 1
.IC V(W_3_26_2) = 1 V(W_3_26_2_bar) = 0
.IC V(W_3_26_3) = 0 V(W_3_26_3_bar) = 1
.IC V(W_3_26_4) = 1 V(W_3_26_4_bar) = 0
.IC V(W_3_27_1) = 0 V(W_3_27_1_bar) = 1
.IC V(W_3_27_2) = 1 V(W_3_27_2_bar) = 0
.IC V(W_3_27_3) = 0 V(W_3_27_3_bar) = 1
.IC V(W_3_27_4) = 1 V(W_3_27_4_bar) = 0
.IC V(W_3_28_1) = 0 V(W_3_28_1_bar) = 1
.IC V(W_3_28_2) = 1 V(W_3_28_2_bar) = 0
.IC V(W_3_28_3) = 0 V(W_3_28_3_bar) = 1
.IC V(W_3_28_4) = 1 V(W_3_28_4_bar) = 0
.IC V(W_3_29_1) = 0 V(W_3_29_1_bar) = 1
.IC V(W_3_29_2) = 1 V(W_3_29_2_bar) = 0
.IC V(W_3_29_3) = 0 V(W_3_29_3_bar) = 1
.IC V(W_3_29_4) = 1 V(W_3_29_4_bar) = 0
.IC V(W_3_30_1) = 0 V(W_3_30_1_bar) = 1
.IC V(W_3_30_2) = 1 V(W_3_30_2_bar) = 0
.IC V(W_3_30_3) = 0 V(W_3_30_3_bar) = 1
.IC V(W_3_30_4) = 1 V(W_3_30_4_bar) = 0
.IC V(W_3_31_1) = 0 V(W_3_31_1_bar) = 1
.IC V(W_3_31_2) = 1 V(W_3_31_2_bar) = 0
.IC V(W_3_31_3) = 0 V(W_3_31_3_bar) = 1
.IC V(W_3_31_4) = 1 V(W_3_31_4_bar) = 0
.IC V(W_3_32_1) = 0 V(W_3_32_1_bar) = 1
.IC V(W_3_32_2) = 1 V(W_3_32_2_bar) = 0
.IC V(W_3_32_3) = 0 V(W_3_32_3_bar) = 1
.IC V(W_3_32_4) = 1 V(W_3_32_4_bar) = 0
.IC V(W_4_1_1) = 0 V(W_4_1_1_bar) = 1
.IC V(W_4_1_2) = 1 V(W_4_1_2_bar) = 0
.IC V(W_4_1_3) = 0 V(W_4_1_3_bar) = 1
.IC V(W_4_1_4) = 1 V(W_4_1_4_bar) = 0
.IC V(W_4_2_1) = 0 V(W_4_2_1_bar) = 1
.IC V(W_4_2_2) = 1 V(W_4_2_2_bar) = 0
.IC V(W_4_2_3) = 0 V(W_4_2_3_bar) = 1
.IC V(W_4_2_4) = 1 V(W_4_2_4_bar) = 0
.IC V(W_4_3_1) = 0 V(W_4_3_1_bar) = 1
.IC V(W_4_3_2) = 1 V(W_4_3_2_bar) = 0
.IC V(W_4_3_3) = 0 V(W_4_3_3_bar) = 1
.IC V(W_4_3_4) = 1 V(W_4_3_4_bar) = 0
.IC V(W_4_4_1) = 0 V(W_4_4_1_bar) = 1
.IC V(W_4_4_2) = 1 V(W_4_4_2_bar) = 0
.IC V(W_4_4_3) = 0 V(W_4_4_3_bar) = 1
.IC V(W_4_4_4) = 1 V(W_4_4_4_bar) = 0
.IC V(W_4_5_1) = 0 V(W_4_5_1_bar) = 1
.IC V(W_4_5_2) = 1 V(W_4_5_2_bar) = 0
.IC V(W_4_5_3) = 0 V(W_4_5_3_bar) = 1
.IC V(W_4_5_4) = 1 V(W_4_5_4_bar) = 0
.IC V(W_4_6_1) = 0 V(W_4_6_1_bar) = 1
.IC V(W_4_6_2) = 1 V(W_4_6_2_bar) = 0
.IC V(W_4_6_3) = 0 V(W_4_6_3_bar) = 1
.IC V(W_4_6_4) = 1 V(W_4_6_4_bar) = 0
.IC V(W_4_7_1) = 0 V(W_4_7_1_bar) = 1
.IC V(W_4_7_2) = 1 V(W_4_7_2_bar) = 0
.IC V(W_4_7_3) = 0 V(W_4_7_3_bar) = 1
.IC V(W_4_7_4) = 1 V(W_4_7_4_bar) = 0
.IC V(W_4_8_1) = 0 V(W_4_8_1_bar) = 1
.IC V(W_4_8_2) = 1 V(W_4_8_2_bar) = 0
.IC V(W_4_8_3) = 0 V(W_4_8_3_bar) = 1
.IC V(W_4_8_4) = 1 V(W_4_8_4_bar) = 0
.IC V(W_4_9_1) = 0 V(W_4_9_1_bar) = 1
.IC V(W_4_9_2) = 1 V(W_4_9_2_bar) = 0
.IC V(W_4_9_3) = 0 V(W_4_9_3_bar) = 1
.IC V(W_4_9_4) = 1 V(W_4_9_4_bar) = 0
.IC V(W_4_10_1) = 0 V(W_4_10_1_bar) = 1
.IC V(W_4_10_2) = 1 V(W_4_10_2_bar) = 0
.IC V(W_4_10_3) = 0 V(W_4_10_3_bar) = 1
.IC V(W_4_10_4) = 1 V(W_4_10_4_bar) = 0
.IC V(W_4_11_1) = 0 V(W_4_11_1_bar) = 1
.IC V(W_4_11_2) = 1 V(W_4_11_2_bar) = 0
.IC V(W_4_11_3) = 0 V(W_4_11_3_bar) = 1
.IC V(W_4_11_4) = 1 V(W_4_11_4_bar) = 0
.IC V(W_4_12_1) = 0 V(W_4_12_1_bar) = 1
.IC V(W_4_12_2) = 1 V(W_4_12_2_bar) = 0
.IC V(W_4_12_3) = 0 V(W_4_12_3_bar) = 1
.IC V(W_4_12_4) = 1 V(W_4_12_4_bar) = 0
.IC V(W_4_13_1) = 0 V(W_4_13_1_bar) = 1
.IC V(W_4_13_2) = 1 V(W_4_13_2_bar) = 0
.IC V(W_4_13_3) = 0 V(W_4_13_3_bar) = 1
.IC V(W_4_13_4) = 1 V(W_4_13_4_bar) = 0
.IC V(W_4_14_1) = 0 V(W_4_14_1_bar) = 1
.IC V(W_4_14_2) = 1 V(W_4_14_2_bar) = 0
.IC V(W_4_14_3) = 0 V(W_4_14_3_bar) = 1
.IC V(W_4_14_4) = 1 V(W_4_14_4_bar) = 0
.IC V(W_4_15_1) = 0 V(W_4_15_1_bar) = 1
.IC V(W_4_15_2) = 1 V(W_4_15_2_bar) = 0
.IC V(W_4_15_3) = 0 V(W_4_15_3_bar) = 1
.IC V(W_4_15_4) = 1 V(W_4_15_4_bar) = 0
.IC V(W_4_16_1) = 0 V(W_4_16_1_bar) = 1
.IC V(W_4_16_2) = 1 V(W_4_16_2_bar) = 0
.IC V(W_4_16_3) = 0 V(W_4_16_3_bar) = 1
.IC V(W_4_16_4) = 1 V(W_4_16_4_bar) = 0
.IC V(W_4_17_1) = 0 V(W_4_17_1_bar) = 1
.IC V(W_4_17_2) = 1 V(W_4_17_2_bar) = 0
.IC V(W_4_17_3) = 0 V(W_4_17_3_bar) = 1
.IC V(W_4_17_4) = 1 V(W_4_17_4_bar) = 0
.IC V(W_4_18_1) = 0 V(W_4_18_1_bar) = 1
.IC V(W_4_18_2) = 1 V(W_4_18_2_bar) = 0
.IC V(W_4_18_3) = 0 V(W_4_18_3_bar) = 1
.IC V(W_4_18_4) = 1 V(W_4_18_4_bar) = 0
.IC V(W_4_19_1) = 0 V(W_4_19_1_bar) = 1
.IC V(W_4_19_2) = 1 V(W_4_19_2_bar) = 0
.IC V(W_4_19_3) = 0 V(W_4_19_3_bar) = 1
.IC V(W_4_19_4) = 1 V(W_4_19_4_bar) = 0
.IC V(W_4_20_1) = 0 V(W_4_20_1_bar) = 1
.IC V(W_4_20_2) = 1 V(W_4_20_2_bar) = 0
.IC V(W_4_20_3) = 0 V(W_4_20_3_bar) = 1
.IC V(W_4_20_4) = 1 V(W_4_20_4_bar) = 0
.IC V(W_4_21_1) = 0 V(W_4_21_1_bar) = 1
.IC V(W_4_21_2) = 1 V(W_4_21_2_bar) = 0
.IC V(W_4_21_3) = 0 V(W_4_21_3_bar) = 1
.IC V(W_4_21_4) = 1 V(W_4_21_4_bar) = 0
.IC V(W_4_22_1) = 0 V(W_4_22_1_bar) = 1
.IC V(W_4_22_2) = 1 V(W_4_22_2_bar) = 0
.IC V(W_4_22_3) = 0 V(W_4_22_3_bar) = 1
.IC V(W_4_22_4) = 1 V(W_4_22_4_bar) = 0
.IC V(W_4_23_1) = 0 V(W_4_23_1_bar) = 1
.IC V(W_4_23_2) = 1 V(W_4_23_2_bar) = 0
.IC V(W_4_23_3) = 0 V(W_4_23_3_bar) = 1
.IC V(W_4_23_4) = 1 V(W_4_23_4_bar) = 0
.IC V(W_4_24_1) = 0 V(W_4_24_1_bar) = 1
.IC V(W_4_24_2) = 1 V(W_4_24_2_bar) = 0
.IC V(W_4_24_3) = 0 V(W_4_24_3_bar) = 1
.IC V(W_4_24_4) = 1 V(W_4_24_4_bar) = 0
.IC V(W_4_25_1) = 0 V(W_4_25_1_bar) = 1
.IC V(W_4_25_2) = 1 V(W_4_25_2_bar) = 0
.IC V(W_4_25_3) = 0 V(W_4_25_3_bar) = 1
.IC V(W_4_25_4) = 1 V(W_4_25_4_bar) = 0
.IC V(W_4_26_1) = 0 V(W_4_26_1_bar) = 1
.IC V(W_4_26_2) = 1 V(W_4_26_2_bar) = 0
.IC V(W_4_26_3) = 0 V(W_4_26_3_bar) = 1
.IC V(W_4_26_4) = 1 V(W_4_26_4_bar) = 0
.IC V(W_4_27_1) = 0 V(W_4_27_1_bar) = 1
.IC V(W_4_27_2) = 1 V(W_4_27_2_bar) = 0
.IC V(W_4_27_3) = 0 V(W_4_27_3_bar) = 1
.IC V(W_4_27_4) = 1 V(W_4_27_4_bar) = 0
.IC V(W_4_28_1) = 0 V(W_4_28_1_bar) = 1
.IC V(W_4_28_2) = 1 V(W_4_28_2_bar) = 0
.IC V(W_4_28_3) = 0 V(W_4_28_3_bar) = 1
.IC V(W_4_28_4) = 1 V(W_4_28_4_bar) = 0
.IC V(W_4_29_1) = 0 V(W_4_29_1_bar) = 1
.IC V(W_4_29_2) = 1 V(W_4_29_2_bar) = 0
.IC V(W_4_29_3) = 0 V(W_4_29_3_bar) = 1
.IC V(W_4_29_4) = 1 V(W_4_29_4_bar) = 0
.IC V(W_4_30_1) = 0 V(W_4_30_1_bar) = 1
.IC V(W_4_30_2) = 1 V(W_4_30_2_bar) = 0
.IC V(W_4_30_3) = 0 V(W_4_30_3_bar) = 1
.IC V(W_4_30_4) = 1 V(W_4_30_4_bar) = 0
.IC V(W_4_31_1) = 0 V(W_4_31_1_bar) = 1
.IC V(W_4_31_2) = 1 V(W_4_31_2_bar) = 0
.IC V(W_4_31_3) = 0 V(W_4_31_3_bar) = 1
.IC V(W_4_31_4) = 1 V(W_4_31_4_bar) = 0
.IC V(W_4_32_1) = 0 V(W_4_32_1_bar) = 1
.IC V(W_4_32_2) = 1 V(W_4_32_2_bar) = 0
.IC V(W_4_32_3) = 0 V(W_4_32_3_bar) = 1
.IC V(W_4_32_4) = 1 V(W_4_32_4_bar) = 0

.end
